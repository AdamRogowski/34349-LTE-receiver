library IEEE;
  use work.complex_pkg.all;

package input_data is

  constant INPUT_DATA_2048_16QAM_CLEAR : complex_array(0 to 2047) := (
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.637595835525, 0.635642710525),
    to_complex(- 1.269329299991, 1.277141799991),
    to_complex(- 0.213181655259, - 0.211228530259),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.128298020250, 0.126344895250),
    to_complex(- 0.420494947286, 0.428307447286),
    to_complex(- 0.091918748841, - 0.089965623841),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.071707598622, 0.069754473622),
    to_complex(- 0.250721684926, 0.258534184926),
    to_complex(- 0.058845594387, - 0.056892469387),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.049940822593, 0.047987697593),
    to_complex(- 0.177957149482, 0.185769649482),
    to_complex(- 0.043410390253, - 0.041457265253),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.038416295193, 0.036463170193),
    to_complex(- 0.137528856024, 0.145341356024),
    to_complex(- 0.034473378260, - 0.032520253260),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.031281302833, 0.029328177833),
    to_complex(- 0.111798854027, 0.119611354027),
    to_complex(- 0.028644197202, - 0.026691072202),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.026428868603, 0.024475743603),
    to_complex(- 0.093983316292, 0.101795816292),
    to_complex(- 0.024541588793, - 0.022588463793),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.022914485594, 0.020961360594),
    to_complex(- 0.080916456729, 0.088728956729),
    to_complex(- 0.021497202231, - 0.019544077231),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.020251589629, 0.018298464629),
    to_complex(- 0.070922270882, 0.078734770882),
    to_complex(- 0.019148218499, - 0.017195093499),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.018164022645, 0.016210897645),
    to_complex(- 0.063030440328, 0.070842940328),
    to_complex(- 0.017280667393, - 0.015327542393),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.016483395569, 0.014530270569),
    to_complex(- 0.056640291713, 0.064452791713),
    to_complex(- 0.015760195518, - 0.013807070518),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.015101190990, 0.013148065990),
    to_complex(- 0.051360081505, 0.059172581505),
    to_complex(- 0.014498186796, - 0.012545061796),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.013944325739, 0.011991200739),
    to_complex(- 0.046923424060, 0.054735924060),
    to_complex(- 0.013433826260, - 0.011480701260),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.012961779486, 0.011008654486),
    to_complex(- 0.043142862780, 0.050955362780),
    to_complex(- 0.012523990562, - 0.010570865562),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.012116853385, 0.010163728385),
    to_complex(- 0.039882653199, 0.047695153199),
    to_complex(- 0.011737250813, - 0.009784125813),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.011382474511, 0.009429349511),
    to_complex(- 0.037042081647, 0.044854581647),
    to_complex(- 0.011050160057, - 0.009097035057),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.010738234036, 0.008785109036),
    to_complex(- 0.034544849863, 0.042357349863),
    to_complex(- 0.010444870603, - 0.008491745603),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.010168455605, 0.008215330605),
    to_complex(- 0.032332099158, 0.040144599158),
    to_complex(- 0.009907556767, - 0.007954431767),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.009660898773, 0.007707773773),
    to_complex(- 0.030357697021, 0.038170197021),
    to_complex(- 0.009427342340, - 0.007474217340),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.009205866554, 0.007252741554),
    to_complex(- 0.028584973994, 0.036397473994),
    to_complex(- 0.008995553882, - 0.007042428882),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.008795577413, 0.006842452413),
    to_complex(- 0.026984415612, 0.034796915612),
    to_complex(- 0.008605189936, - 0.006652064936),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.008423714566, 0.006470589566),
    to_complex(- 0.025531998452, 0.033344498452),
    to_complex(- 0.008250536662, - 0.006297411662),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.008085096829, 0.006131971829),
    to_complex(- 0.024207969896, 0.032020469896),
    to_complex(- 0.007926884849, - 0.005973759849),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.007775434394, 0.005822309394),
    to_complex(- 0.022995939456, 0.030808439456),
    to_complex(- 0.007630318408, - 0.005677193408),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.007491145051, 0.005538020051),
    to_complex(- 0.021882192621, 0.029694692621),
    to_complex(- 0.007357554149, - 0.005404429149),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.007229214058, 0.005276089058),
    to_complex(- 0.020855166156, 0.028667666156),
    to_complex(- 0.007105818889, - 0.005152693889),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.006987086062, 0.005033961062),
    to_complex(- 0.019905042202, 0.027717542202),
    to_complex(- 0.006872754121, - 0.004919629121),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.006762580801, 0.004809455801),
    to_complex(- 0.019023430933, 0.026835930933),
    to_complex(- 0.006656341296, - 0.004703216296),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.006553826718, 0.004600701718),
    to_complex(- 0.018203120025, 0.026015620025),
    to_complex(- 0.006454842707, - 0.004501717707),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.006359208193, 0.004406083193),
    to_complex(- 0.017437875081, 0.025250375081),
    to_complex(- 0.006266754280, - 0.004313629280),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.006177323236, 0.004224198236),
    to_complex(- 0.016722279311, 0.024534779311),
    to_complex(- 0.006090767590, - 0.004137642590),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.006006949308, 0.004053824308),
    to_complex(- 0.016051603757, 0.023864103757),
    to_complex(- 0.005925739051, - 0.003972614051),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.005847015499, 0.003893890499),
    to_complex(- 0.015421701470, 0.023234201470),
    to_complex(- 0.005770664744, - 0.003817539744),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.005696579726, 0.003743454726),
    to_complex(- 0.014828920645, 0.022641420645),
    to_complex(- 0.005624659732, - 0.003671534732),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.005554809928, 0.003601684928),
    to_complex(- 0.014270032858, 0.022082532858),
    to_complex(- 0.005486940938, - 0.003533815938),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.005420968456, 0.003467843456),
    to_complex(- 0.013742173440, 0.021554673440),
    to_complex(- 0.005356812895, - 0.003403687895),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.005294399056, 0.003341274056),
    to_complex(- 0.013242791641, 0.021055291641),
    to_complex(- 0.005233655834, - 0.003280530834),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.005174515940, 0.003221390940),
    to_complex(- 0.012769608778, 0.020582108778),
    to_complex(- 0.005116915650, - 0.003163790650),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.005060794574, 0.003107669574),
    to_complex(- 0.012320582903, 0.020133082903),
    to_complex(- 0.005006095435, - 0.003052970435),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.004952763878, 0.002999638878),
    to_complex(- 0.011893878832, 0.019706378832),
    to_complex(- 0.004900748279, - 0.002947623279),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.004849999583, 0.002896874583),
    to_complex(- 0.011487842622, 0.019300342622),
    to_complex(- 0.004800471139, - 0.002847346139),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.004752118560, 0.002798993560),
    to_complex(- 0.011100979732, 0.018913479732),
    to_complex(- 0.004704899583, - 0.002751774583),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.004658773947, 0.002705648947),
    to_complex(- 0.010731936275, 0.018544436275),
    to_complex(- 0.004613703275, - 0.002660578275),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.004569650961, 0.002616525961),
    to_complex(- 0.010379482843, 0.018191982843),
    to_complex(- 0.004526582077, - 0.002573457077),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.004484463269, 0.002531338269),
    to_complex(- 0.010042500528, 0.017855000528),
    to_complex(- 0.004443262678, - 0.002490137678),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.004402949848, 0.002449824848),
    to_complex(- 0.009719968773, 0.017532468773),
    to_complex(- 0.004363495658, - 0.002410370658),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.004324872245, 0.002371747245),
    to_complex(- 0.009410954802, 0.017223454802),
    to_complex(- 0.004287052938, - 0.002333927938),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.004250012193, 0.002296887193),
    to_complex(- 0.009114604375, 0.016927104375),
    to_complex(- 0.004213725538, - 0.002260600538),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.004178169515, 0.002225044515),
    to_complex(- 0.008830133696, 0.016642633696),
    to_complex(- 0.004143321627, - 0.002190196627),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.004109160291, 0.002156035291),
    to_complex(- 0.008556822293, 0.016369322293),
    to_complex(- 0.004075664791, - 0.002122539791),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.004042815236, 0.002089690236),
    to_complex(- 0.008294006750, 0.016106506750),
    to_complex(- 0.004010592519, - 0.002057467519),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.003978978278, 0.002025853278),
    to_complex(- 0.008041075171, 0.015853575171),
    to_complex(- 0.003947954860, - 0.001994829860),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.003917505289, 0.001964380289),
    to_complex(- 0.007797462267, 0.015609962267),
    to_complex(- 0.003887613230, - 0.001934488230),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.003858262964, 0.001905137964),
    to_complex(- 0.007562645004, 0.015375145004),
    to_complex(- 0.003829439355, - 0.001876314355),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.003801127826, 0.001848002826),
    to_complex(- 0.007336138727, 0.015148638727),
    to_complex(- 0.003773314331, - 0.001820189331),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.003745985334, 0.001792860334),
    to_complex(- 0.007117493699, 0.014929993699),
    to_complex(- 0.003719127783, - 0.001766002783),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.003692729090, 0.001739604090),
    to_complex(- 0.006906292015, 0.014718792015),
    to_complex(- 0.003666777112, - 0.001713652112),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.003641260127, 0.001688135127),
    to_complex(- 0.006702144829, 0.014514644829),
    to_complex(- 0.003616166823, - 0.001663041823),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.003591486273, 0.001638361273),
    to_complex(- 0.006504689876, 0.014317189876),
    to_complex(- 0.003567207923, - 0.001614082923),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.003543321575, 0.001590196575),
    to_complex(- 0.006313589233, 0.014126089233),
    to_complex(- 0.003519817372, - 0.001566692372),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.003496685783, 0.001543560783),
    to_complex(- 0.006128527311, 0.013941027311),
    to_complex(- 0.003473917594, - 0.001520792594),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.003451503888, 0.001498378888),
    to_complex(- 0.005949209038, 0.013761709038),
    to_complex(- 0.003429436039, - 0.001476311039),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.003407705696, 0.001454580696),
    to_complex(- 0.005775358215, 0.013587858215),
    to_complex(- 0.003386304777, - 0.001433179777),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.003365225452, 0.001412100452),
    to_complex(- 0.005606716035, 0.013419216035),
    to_complex(- 0.003344460139, - 0.001391335139),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.003324001491, 0.001370876491),
    to_complex(- 0.005443039729, 0.013255539729),
    to_complex(- 0.003303842387, - 0.001350717387),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.003283975926, 0.001330850926),
    to_complex(- 0.005284101347, 0.013096601347),
    to_complex(- 0.003264395415, - 0.001311270415),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.003245094363, 0.001291969363),
    to_complex(- 0.005129686641, 0.012942186641),
    to_complex(- 0.003226066476, - 0.001272941476),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.003207305643, 0.001254180643),
    to_complex(- 0.004979594048, 0.012792094048),
    to_complex(- 0.003188805936, - 0.001235680936),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.003170561599, 0.001217436599),
    to_complex(- 0.004833633770, 0.012646133770),
    to_complex(- 0.003152567046, - 0.001199442046),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.003134816848, 0.001181691848),
    to_complex(- 0.004691626920, 0.012504126920),
    to_complex(- 0.003117305736, - 0.001164180736),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.003100028587, 0.001146903587),
    to_complex(- 0.004553404754, 0.012365904754),
    to_complex(- 0.003082980426, - 0.001129855426),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.003066156414, 0.001113031414),
    to_complex(- 0.004418807960, 0.012231307960),
    to_complex(- 0.003049551850, - 0.001096426850),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.003033162162, 0.001080037162),
    to_complex(- 0.004287686005, 0.012100186005),
    to_complex(- 0.003016982902, - 0.001063857902),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.003001009745, 0.001047884745),
    to_complex(- 0.004159896542, 0.011972396542),
    to_complex(- 0.002985238483, - 0.001032113483),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.002969665021, 0.001016540021),
    to_complex(- 0.004035304858, 0.011847804858),
    to_complex(- 0.002954285372, - 0.001001160372),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.002939095658, 0.000985970658),
    to_complex(- 0.003913783367, 0.011726283367),
    to_complex(- 0.002924092100, - 0.000970967100),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.002909271021, 0.000956146021),
    to_complex(- 0.003795211147, 0.011607711147),
    to_complex(- 0.002894628836, - 0.000941503836),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.002880162056, 0.000927037056),
    to_complex(- 0.003679473509, 0.011491973509),
    to_complex(- 0.002865867281, - 0.000912742281),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.002851741196, 0.000898616196),
    to_complex(- 0.003566461600, 0.011378961600),
    to_complex(- 0.002837780572, - 0.000884655572),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.002823982260, 0.000870857260),
    to_complex(- 0.003456072034, 0.011268572034),
    to_complex(- 0.002810343190, - 0.000857218190),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.002796860370, 0.000843735370),
    to_complex(- 0.003348206556, 0.011160706556),
    to_complex(- 0.002783530881, - 0.000830405881),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.002770351874, 0.000817226874),
    to_complex(- 0.003242771724, 0.011055271724),
    to_complex(- 0.002757320572, - 0.000804195572),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.002744434265, 0.000791309265),
    to_complex(- 0.003139678618, 0.010952178618),
    to_complex(- 0.002731690306, - 0.000778565306),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.002719086115, 0.000765961115),
    to_complex(- 0.003038842571, 0.010851342571),
    to_complex(- 0.002706619172, - 0.000753494172),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.002694287015, 0.000741162015),
    to_complex(- 0.002940182915, 0.010752682915),
    to_complex(- 0.002682087243, - 0.000728962243),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.002670017508, 0.000716892508),
    to_complex(- 0.002843622748, 0.010656122748),
    to_complex(- 0.002658075520, - 0.000704950520),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.002646259040, 0.000693134040),
    to_complex(- 0.002749088717, 0.010561588717),
    to_complex(- 0.002634565879, - 0.000681440879),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.002622993902, 0.000669868902),
    to_complex(- 0.002656510811, 0.010469010811),
    to_complex(- 0.002611541020, - 0.000658416020),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.002600205190, 0.000647080190),
    to_complex(- 0.002565822181, 0.010378322181),
    to_complex(- 0.002588984419, - 0.000635859419),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.002577876754, 0.000624751754),
    to_complex(- 0.002476958953, 0.010289458953),
    to_complex(- 0.002566880288, - 0.000613755288),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.002555993155, 0.000602868155),
    to_complex(- 0.002389860070, 0.010202360070),
    to_complex(- 0.002545213532, - 0.000592088532),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.002534539634, 0.000581414634),
    to_complex(- 0.002304467136, 0.010116967136),
    to_complex(- 0.002523969714, - 0.000570844714),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.002513502065, 0.000560377065),
    to_complex(- 0.002220724273, 0.010033224273),
    to_complex(- 0.002503135015, - 0.000550010015),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.002492866930, 0.000539741930),
    to_complex(- 0.002138577986, 0.009951077986),
    to_complex(- 0.002482696207, - 0.000529571207),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.002472621279, 0.000519496279),
    to_complex(- 0.002057977034, 0.009870477034),
    to_complex(- 0.002462640614, - 0.000509515614),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.002452752708, 0.000499627708),
    to_complex(- 0.001978872317, 0.009791372317),
    to_complex(- 0.002442956091, - 0.000489831091),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.002433249323, 0.000480124323),
    to_complex(- 0.001901216762, 0.009713716762),
    to_complex(- 0.002423630993, - 0.000470505993),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.002414099720, 0.000460974720),
    to_complex(- 0.001824965219, 0.009637465219),
    to_complex(- 0.002404654149, - 0.000451529149),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.002395292954, 0.000442167954),
    to_complex(- 0.001750074363, 0.009562574363),
    to_complex(- 0.002386014836, - 0.000432889836),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.002376818523, 0.000423693523),
    to_complex(- 0.001676502604, 0.009489002604),
    to_complex(- 0.002367702764, - 0.000414577764),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.002358666339, 0.000405541339),
    to_complex(- 0.001604209999, 0.009416709999),
    to_complex(- 0.002349708046, - 0.000396583046),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.002340826712, 0.000387701712),
    to_complex(- 0.001533158172, 0.009345658172),
    to_complex(- 0.002332021183, - 0.000378896183),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.002323290330, 0.000370165330),
    to_complex(- 0.001463310237, 0.009275810237),
    to_complex(- 0.002314633044, - 0.000361508044),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.002306048238, 0.000352923238),
    to_complex(- 0.001394630723, 0.009207130723),
    to_complex(- 0.002297534846, - 0.000344409846),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.002289091823, 0.000335966823),
    to_complex(- 0.001327085514, 0.009139585514),
    to_complex(- 0.002280718143, - 0.000327593143),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.002272412799, 0.000319287799),
    to_complex(- 0.001260641774, 0.009073141774),
    to_complex(- 0.002264174804, - 0.000311049804),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.002256003188, 0.000302878188),
    to_complex(- 0.001195267898, 0.009007767898),
    to_complex(- 0.002247897001, - 0.000294772001),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.002239855309, 0.000286730309),
    to_complex(- 0.001130933446, 0.008943433446),
    to_complex(- 0.002231877196, - 0.000278752196),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.002223961762, 0.000270836762),
    to_complex(- 0.001067609092, 0.008880109092),
    to_complex(- 0.002216108124, - 0.000262983124),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.002208315416, 0.000255190416),
    to_complex(- 0.001005266576, 0.008817766576),
    to_complex(- 0.002200582786, - 0.000247457786),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.002192909398, 0.000239784398),
    to_complex(- 0.000943878651, 0.008756378651),
    to_complex(- 0.002185294431, - 0.000232169431),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.002177737079, 0.000224612079),
    to_complex(- 0.000883419041, 0.008695919041),
    to_complex(- 0.002170236549, - 0.000217111549),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.002162792064, 0.000209667064),
    to_complex(- 0.000823862396, 0.008636362396),
    to_complex(- 0.002155402859, - 0.000202277859),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.002148068183, 0.000194943183),
    to_complex(- 0.000765184251, 0.008577684251),
    to_complex(- 0.002140787299, - 0.000187662299),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.002133559480, 0.000180434480),
    to_complex(- 0.000707360990, 0.008519860990),
    to_complex(- 0.002126384015, - 0.000173259015),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.002119260203, 0.000166135203),
    to_complex(- 0.000650369804, 0.008462869804),
    to_complex(- 0.002112187355, - 0.000159062355),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.002105164796, 0.000152039796),
    to_complex(- 0.000594188662, 0.008406688662),
    to_complex(- 0.002098191859, - 0.000145066859),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.002091267891, 0.000138142891),
    to_complex(- 0.000538796274, 0.008351296274),
    to_complex(- 0.002084392248, - 0.000131267248),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.002077564299, 0.000124439299),
    to_complex(- 0.000484172060, 0.008296672060),
    to_complex(- 0.002070783422, - 0.000117658422),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.002064049005, 0.000110924005),
    to_complex(- 0.000430296122, 0.008242796122),
    to_complex(- 0.002057360447, - 0.000104235447),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.002050717156, 0.000097592156),
    to_complex(- 0.000377149215, 0.008189649215),
    to_complex(- 0.002044118551, - 0.000090993551),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.002037564059, 0.000084439059),
    to_complex(- 0.000324712718, 0.008137212718),
    to_complex(- 0.002031053118, - 0.000077928118),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.002024585173, 0.000071460173),
    to_complex(- 0.000272968613, 0.008085468613),
    to_complex(- 0.002018159679, - 0.000065034679),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.002011776100, 0.000058651100),
    to_complex(- 0.000221899454, 0.008034399454),
    to_complex(- 0.002005433908, - 0.000052308908),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001999132584, 0.000046007584),
    to_complex(- 0.000171488351, 0.007983988351),
    to_complex(- 0.001992871617, - 0.000039746617),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001986650503, 0.000033525503),
    to_complex(- 0.000121718942, 0.007934218942),
    to_complex(- 0.001980468746, - 0.000027343746),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001974325860, 0.000021200860),
    to_complex(- 0.000072575374, 0.007885075374),
    to_complex(- 0.001968221365, - 0.000015096365),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001962154787, 0.000009029787),
    to_complex(- 0.000024042286, 0.007836542286),
    to_complex(- 0.001956125662, - 0.000003000662),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001950133530, - 0.000002991470),
    to_complex(0.000023895215, 0.007788604785),
    to_complex(- 0.001944177942, 0.000008947058),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001938258452, - 0.000014866548),
    to_complex(0.000071251570, 0.007741248430),
    to_complex(- 0.001932374624, 0.000020750376),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001926526025, - 0.000026598975),
    to_complex(0.000118040785, 0.007694459215),
    to_complex(- 0.001920712231, 0.000032412769),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001914932825, - 0.000038192175),
    to_complex(0.000164276448, 0.007648223552),
    to_complex(- 0.001909187394, 0.000043937606),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001903475532, - 0.000049649468),
    to_complex(0.000209971745, 0.007602528255),
    to_complex(- 0.001897796839, 0.000055328161),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001892150921, - 0.000060974079),
    to_complex(0.000255139475, 0.007557360525),
    to_complex(- 0.001886537390, 0.000066587610),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001880955863, - 0.000072169137),
    to_complex(0.000299792066, 0.007512707934),
    to_complex(- 0.001875405964, 0.000077719036),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001869887319, - 0.000083237681),
    to_complex(0.000343941586, 0.007468558414),
    to_complex(- 0.001864399564, 0.000088725436),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001858942337, - 0.000094182663),
    to_complex(0.000387599758, 0.007424900242),
    to_complex(- 0.001853515283, 0.000099609717),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001848118049, - 0.000105006951),
    to_complex(0.000430777971, 0.007381722029),
    to_complex(- 0.001842750291, 0.000110374709),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001837411667, - 0.000115713333),
    to_complex(0.000473487297, 0.007339012703),
    to_complex(- 0.001832101842, 0.000121023158),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001826820483, - 0.000126304517),
    to_complex(0.000515738495, 0.007296761505),
    to_complex(- 0.001821567264, 0.000131557736),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001816341862, - 0.000136783138),
    to_complex(0.000557542028, 0.007254957972),
    to_complex(- 0.001811143959, 0.000141981041),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001805973242, - 0.000147151758),
    to_complex(0.000598908073, 0.007213591927),
    to_complex(- 0.001800829402, 0.000152295598),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001795712133, - 0.000157412867),
    to_complex(0.000639846527, 0.007172653473),
    to_complex(- 0.001790621134, 0.000162503866),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001785556109, - 0.000167568891),
    to_complex(0.000680367022, 0.007132132978),
    to_complex(- 0.001780516764, 0.000172608236),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001775502811, - 0.000177622189),
    to_complex(0.000720478930, 0.007092021070),
    to_complex(- 0.001770513965, 0.000182611035),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001765549944, - 0.000187575056),
    to_complex(0.000760191377, 0.007052308623),
    to_complex(- 0.001760610470, 0.000192514530),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001755695270, - 0.000197429730),
    to_complex(0.000799513246, 0.007012986754),
    to_complex(- 0.001750804074, 0.000202320926),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001745936614, - 0.000207188386),
    to_complex(0.000838453189, 0.006974046811),
    to_complex(- 0.001741092627, 0.000212032373),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001736271854, - 0.000216853146),
    to_complex(0.000877019632, 0.006935480368),
    to_complex(- 0.001731474037, 0.000221650963),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001726698924, - 0.000226426076),
    to_complex(0.000915220787, 0.006897279213),
    to_complex(- 0.001721946264, 0.000231178736),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001717215811, - 0.000235909189),
    to_complex(0.000953064656, 0.006859435344),
    to_complex(- 0.001712507321, 0.000240617679),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001707820553, - 0.000245304447),
    to_complex(0.000990559037, 0.006821940963),
    to_complex(- 0.001703155270, 0.000249969730),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001698511237, - 0.000254613763),
    to_complex(0.001027711535, 0.006784788465),
    to_complex(- 0.001693888222, 0.000259236778),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001689285997, - 0.000263839003),
    to_complex(0.001064529563, 0.006747970437),
    to_complex(- 0.001684704335, 0.000268420665),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001680143014, - 0.000272981986),
    to_complex(0.001101020354, 0.006711479646),
    to_complex(- 0.001675601812, 0.000277523188),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001671080513, - 0.000282044487),
    to_complex(0.001137190962, 0.006675309038),
    to_complex(- 0.001666578901, 0.000286546099),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001662096763, - 0.000291028237),
    to_complex(0.001173048272, 0.006639451728),
    to_complex(- 0.001657633891, 0.000295491109),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001653190075, - 0.000299934925),
    to_complex(0.001208599002, 0.006603900998),
    to_complex(- 0.001648765112, 0.000304359888),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001644358798, - 0.000308766202),
    to_complex(0.001243849710, 0.006568650290),
    to_complex(- 0.001639970935, 0.000313154065),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001635601323, - 0.000317523677),
    to_complex(0.001278806799, 0.006533693201),
    to_complex(- 0.001631249768, 0.000321875232),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001626916076, - 0.000326208924),
    to_complex(0.001313476521, 0.006499023479),
    to_complex(- 0.001622600057, 0.000330524943),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001618301523, - 0.000334823477),
    to_complex(0.001347864986, 0.006464635014),
    to_complex(- 0.001614020285, 0.000339104715),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001609756162, - 0.000343368838),
    to_complex(0.001381978160, 0.006430521840),
    to_complex(- 0.001605508969, 0.000347616031),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001601278527, - 0.000351846473),
    to_complex(0.001415821873, 0.006396678127),
    to_complex(- 0.001597064658, 0.000356060342),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001592867186, - 0.000360257814),
    to_complex(0.001449401825, 0.006363098175),
    to_complex(- 0.001588685936, 0.000364439064),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001584520737, - 0.000368604263),
    to_complex(0.001482723586, 0.006329776414),
    to_complex(- 0.001580371419, 0.000372753581),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001576237813, - 0.000376887187),
    to_complex(0.001515792602, 0.006296707398),
    to_complex(- 0.001572119752, 0.000381005248),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001568017072, - 0.000385107928),
    to_complex(0.001548614202, 0.006263885798),
    to_complex(- 0.001563929611, 0.000389195389),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001559857207, - 0.000393267793),
    to_complex(0.001581193595, 0.006231306405),
    to_complex(- 0.001555799701, 0.000397325299),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001551756935, - 0.000401368065),
    to_complex(0.001613535878, 0.006198964122),
    to_complex(- 0.001547728753, 0.000405396247),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001543715002, - 0.000409409998),
    to_complex(0.001645646040, 0.006166853960),
    to_complex(- 0.001539715528, 0.000413409472),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001535730182, - 0.000417394818),
    to_complex(0.001677528964, 0.006134971036),
    to_complex(- 0.001531758812, 0.000421366188),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001527801273, - 0.000425323727),
    to_complex(0.001709189427, 0.006103310573),
    to_complex(- 0.001523857416, 0.000429267584),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001519927099, - 0.000433197901),
    to_complex(0.001740632111, 0.006071867889),
    to_complex(- 0.001516010177, 0.000437114823),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001512106509, - 0.000441018491),
    to_complex(0.001771861597, 0.006040638403),
    to_complex(- 0.001508215954, 0.000444909046),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001504338374, - 0.000448786626),
    to_complex(0.001802882374, 0.006009617626),
    to_complex(- 0.001500473631, 0.000452651369),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001496621590, - 0.000456503410),
    to_complex(0.001833698841, 0.005978801159),
    to_complex(- 0.001492782115, 0.000460342885),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001488955073, - 0.000464169927),
    to_complex(0.001864315308, 0.005948184692),
    to_complex(- 0.001485140332, 0.000467984668),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001481337762, - 0.000471787238),
    to_complex(0.001894735997, 0.005917764003),
    to_complex(- 0.001477547233, 0.000475577767),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001473768618, - 0.000479356382),
    to_complex(0.001924965050, 0.005887534950),
    to_complex(- 0.001470001788, 0.000483123212),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001466246619, - 0.000486878381),
    to_complex(0.001955006527, 0.005857493473),
    to_complex(- 0.001462502986, 0.000490622014),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001458770766, - 0.000494354234),
    to_complex(0.001984864410, 0.005827635590),
    to_complex(- 0.001455049837, 0.000498075163),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001451340077, - 0.000501784923),
    to_complex(0.002014542605, 0.005797957395),
    to_complex(- 0.001447641368, 0.000505483632),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001443953590, - 0.000509171410),
    to_complex(0.002044044943, 0.005768455057),
    to_complex(- 0.001440276627, 0.000512848373),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001436610361, - 0.000516514639),
    to_complex(0.002073375186, 0.005739124814),
    to_complex(- 0.001432954677, 0.000520170323),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001429309462, - 0.000523815538),
    to_complex(0.002102537023, 0.005709962977),
    to_complex(- 0.001425674601, 0.000527450399),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001422049983, - 0.000531075017),
    to_complex(0.002131534078, 0.005680965922),
    to_complex(- 0.001418435497, 0.000534689503),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001414831031, - 0.000538293969),
    to_complex(0.002160369910, 0.005652130090),
    to_complex(- 0.001411236478, 0.000541888522),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001407651729, - 0.000545473271),
    to_complex(0.002189048012, 0.005623451988),
    to_complex(- 0.001404076676, 0.000549048324),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001400511213, - 0.000552613787),
    to_complex(0.002217571818, 0.005594928182),
    to_complex(- 0.001396955236, 0.000556169764),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001393408639, - 0.000559716361),
    to_complex(0.002245944699, 0.005566555301),
    to_complex(- 0.001389871318, 0.000563253682),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001386343172, - 0.000566781828),
    to_complex(0.002274169970, 0.005538330030),
    to_complex(- 0.001382824098, 0.000570300902),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001379313996, - 0.000573811004),
    to_complex(0.002302250889, 0.005510249111),
    to_complex(- 0.001375812765, 0.000577312235),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001372320306, - 0.000580804694),
    to_complex(0.002330190659, 0.005482309341),
    to_complex(- 0.001368836521, 0.000584288479),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001365361311, - 0.000587763689),
    to_complex(0.002357992430, 0.005454507570),
    to_complex(- 0.001361894581, 0.000591230419),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001358436235, - 0.000594688765),
    to_complex(0.002385659299, 0.005426840701),
    to_complex(- 0.001354986176, 0.000598138824),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001351544311, - 0.000601580689),
    to_complex(0.002413194315, 0.005399305685),
    to_complex(- 0.001348110545, 0.000605014455),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001344684786, - 0.000608440214),
    to_complex(0.002440600477, 0.005371899523),
    to_complex(- 0.001341266942, 0.000611858058),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001337856921, - 0.000615268079),
    to_complex(0.002467880736, 0.005344619264),
    to_complex(- 0.001334454633, 0.000618670367),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001331059986, - 0.000622065014),
    to_complex(0.002495037998, 0.005317462002),
    to_complex(- 0.001327672892, 0.000625452108),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001324293262, - 0.000628831738),
    to_complex(0.002522075124, 0.005290424876),
    to_complex(- 0.001320921008, 0.000632203992),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001317556043, - 0.000635568957),
    to_complex(0.002548994933, 0.005263505067),
    to_complex(- 0.001314198280, 0.000638926720),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001310847632, - 0.000642277368),
    to_complex(0.002575800200, 0.005236699800),
    to_complex(- 0.001307504015, 0.000645620985),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001304167343, - 0.000648957657),
    to_complex(0.002602493661, 0.005210006339),
    to_complex(- 0.001300837532, 0.000652287468),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001297514499, - 0.000655610501),
    to_complex(0.002629078010, 0.005183421990),
    to_complex(- 0.001294198160, 0.000658926840),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001290888433, - 0.000662236567),
    to_complex(0.002655555906, 0.005156944094),
    to_complex(- 0.001287585236, 0.000665539764),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001284288489, - 0.000668836511),
    to_complex(0.002681929968, 0.005130570032),
    to_complex(- 0.001280998109, 0.000672126891),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001277714017, - 0.000675410983),
    to_complex(0.002708202781, 0.005104297219),
    to_complex(- 0.001274436134, 0.000678688866),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001271164380, - 0.000681960620),
    to_complex(0.002734376894, 0.005078123106),
    to_complex(- 0.001267898676, 0.000685226324),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001264638945, - 0.000688486055),
    to_complex(0.002760454821, 0.005052045179),
    to_complex(- 0.001261385109, 0.000691739891),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001258137090, - 0.000694987910),
    to_complex(0.002786439045, 0.005026060955),
    to_complex(- 0.001254894813, 0.000698230187),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001251658201, - 0.000701466799),
    to_complex(0.002812332016, 0.005000167984),
    to_complex(- 0.001248427179, 0.000704697821),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001245201671, - 0.000707923329),
    to_complex(0.002838136153, 0.004974363847),
    to_complex(- 0.001241981603, 0.000711143397),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001238766901, - 0.000714358099),
    to_complex(0.002863853847, 0.004948646153),
    to_complex(- 0.001235557490, 0.000717567510),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001232353298, - 0.000720771702),
    to_complex(0.002889487457, 0.004923012543),
    to_complex(- 0.001229154251, 0.000723970749),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001225960278, - 0.000727164722),
    to_complex(0.002915039317, 0.004897460683),
    to_complex(- 0.001222771305, 0.000730353695),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001219587262, - 0.000733537738),
    to_complex(0.002940511731, 0.004871988269),
    to_complex(- 0.001216408078, 0.000736716922),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001213233680, - 0.000739891320),
    to_complex(0.002965906980, 0.004846593020),
    to_complex(- 0.001210064000, 0.000743061000),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001206898967, - 0.000746226033),
    to_complex(0.002991227316, 0.004821272684),
    to_complex(- 0.001203738511, 0.000749386489),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001200582563, - 0.000752542437),
    to_complex(0.003016474969, 0.004796025031),
    to_complex(- 0.001197431054, 0.000755693946),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001194283916, - 0.000758841084),
    to_complex(0.003041652144, 0.004770847856),
    to_complex(- 0.001191141079, 0.000761983921),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001188002478, - 0.000765122522),
    to_complex(0.003066761025, 0.004745738975),
    to_complex(- 0.001184868043, 0.000768256957),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001181737708, - 0.000771387292),
    to_complex(0.003091803772, 0.004720696228),
    to_complex(- 0.001178611406, 0.000774513594),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001175489070, - 0.000777635930),
    to_complex(0.003116782524, 0.004695717476),
    to_complex(- 0.001172370635, 0.000780754365),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001169256033, - 0.000783868967),
    to_complex(0.003141699400, 0.004670800600),
    to_complex(- 0.001166145201, 0.000786979799),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001163038071, - 0.000790086929),
    to_complex(0.003166556499, 0.004645943501),
    to_complex(- 0.001159934581, 0.000793190419),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001156834663, - 0.000796290337),
    to_complex(0.003191355901, 0.004621144099),
    to_complex(- 0.001153738255, 0.000799386745),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001150645292, - 0.000802479708),
    to_complex(0.003216099668, 0.004596400332),
    to_complex(- 0.001147555711, 0.000805569289),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001144469447, - 0.000808655553),
    to_complex(0.003240789843, 0.004571710157),
    to_complex(- 0.001141386437, 0.000811738563),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001138306619, - 0.000814818381),
    to_complex(0.003265428455, 0.004547071545),
    to_complex(- 0.001135229928, 0.000817895072),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001132156304, - 0.000820968696),
    to_complex(0.003290017513, 0.004522482487),
    to_complex(- 0.001129085683, 0.000824039317),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001126018003, - 0.000827106997),
    to_complex(0.003314559013, 0.004497940987),
    to_complex(- 0.001122953203, 0.000830171797),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001119891220, - 0.000833233780),
    to_complex(0.003339054936, 0.004473445064),
    to_complex(- 0.001116831993, 0.000836293007),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001113775462, - 0.000839349538),
    to_complex(0.003363507249, 0.004448992751),
    to_complex(- 0.001110721565, 0.000842403435),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001107670240, - 0.000845454760),
    to_complex(0.003387917903, 0.004424582097),
    to_complex(- 0.001104621429, 0.000848503571),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001101575069, - 0.000851549931),
    to_complex(0.003412288839, 0.004400211161),
    to_complex(- 0.001098531102, 0.000854593898),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001095489466, - 0.000857635534),
    to_complex(0.003436621984, 0.004375878016),
    to_complex(- 0.001092450102, 0.000860674898),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001089412951, - 0.000863712049),
    to_complex(0.003460919255, 0.004351580745),
    to_complex(- 0.001086377952, 0.000866747048),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001083345047, - 0.000869779953),
    to_complex(0.003485182556, 0.004327317444),
    to_complex(- 0.001080314176, 0.000872810824),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001077285280, - 0.000875839720),
    to_complex(0.003509413782, 0.004303086218),
    to_complex(- 0.001074258301, 0.000878866699),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001071233179, - 0.000881891821),
    to_complex(0.003533614817, 0.004278885183),
    to_complex(- 0.001068209855, 0.000884915145),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001065188273, - 0.000887936727),
    to_complex(0.003557787537, 0.004254712463),
    to_complex(- 0.001062168372, 0.000890956628),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001059150095, - 0.000893974905),
    to_complex(0.003581933809, 0.004230566191),
    to_complex(- 0.001056133384, 0.000896991616),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001053118181, - 0.000900006819),
    to_complex(0.003606055491, 0.004206444509),
    to_complex(- 0.001050104428, 0.000903020572),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001047092068, - 0.000906032932),
    to_complex(0.003630154434, 0.004182345566),
    to_complex(- 0.001044081042, 0.000909043958),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001041071293, - 0.000912053707),
    to_complex(0.003654232484, 0.004158267516),
    to_complex(- 0.001038062763, 0.000915062237),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001035055396, - 0.000918069604),
    to_complex(0.003678291477, 0.004134208523),
    to_complex(- 0.001032049134, 0.000921075866),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001029043920, - 0.000924081080),
    to_complex(0.003702333246, 0.004110166754),
    to_complex(- 0.001026039697, 0.000927085303),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001023036408, - 0.000930088592),
    to_complex(0.003726359619, 0.004086140381),
    to_complex(- 0.001020033995, 0.000933091005),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001017032402, - 0.000936092598),
    to_complex(0.003750372416, 0.004062127584),
    to_complex(- 0.001014031573, 0.000939093427),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001011031450, - 0.000942093550),
    to_complex(0.003774373458, 0.004038126542),
    to_complex(- 0.001008031977, 0.000945093023),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001005033096, - 0.000948091904),
    to_complex(0.003798364557, 0.004014135443),
    to_complex(- 0.001002034752, 0.000951090248),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000999036888, - 0.000954088112),
    to_complex(0.003822347526, 0.003990152474),
    to_complex(- 0.000996039447, 0.000957085553),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000993042373, - 0.000960082627),
    to_complex(0.003846324175, 0.003966175825),
    to_complex(- 0.000990045610, 0.000963079390),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000987049100, - 0.000966075900),
    to_complex(0.003870296310, 0.003942203690),
    to_complex(- 0.000984052787, 0.000969072213),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000981056616, - 0.000972068384),
    to_complex(0.003894265737, 0.003918234263),
    to_complex(- 0.000978060529, 0.000975064471),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000975064471, - 0.000978060529),
    to_complex(0.003918234263, 0.003894265737),
    to_complex(- 0.000972068384, 0.000981056616),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000969072213, - 0.000984052787),
    to_complex(0.003942203690, 0.003870296310),
    to_complex(- 0.000966075900, 0.000987049100),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000963079390, - 0.000990045610),
    to_complex(0.003966175825, 0.003846324175),
    to_complex(- 0.000960082627, 0.000993042373),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000957085553, - 0.000996039447),
    to_complex(0.003990152474, 0.003822347526),
    to_complex(- 0.000954088112, 0.000999036888),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000951090248, - 0.001002034752),
    to_complex(0.004014135443, 0.003798364557),
    to_complex(- 0.000948091904, 0.001005033096),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000945093023, - 0.001008031977),
    to_complex(0.004038126542, 0.003774373458),
    to_complex(- 0.000942093550, 0.001011031450),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000939093427, - 0.001014031573),
    to_complex(0.004062127584, 0.003750372416),
    to_complex(- 0.000936092598, 0.001017032402),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000933091005, - 0.001020033995),
    to_complex(0.004086140381, 0.003726359619),
    to_complex(- 0.000930088592, 0.001023036408),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000927085303, - 0.001026039697),
    to_complex(0.004110166754, 0.003702333246),
    to_complex(- 0.000924081080, 0.001029043920),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000921075866, - 0.001032049134),
    to_complex(0.004134208523, 0.003678291477),
    to_complex(- 0.000918069604, 0.001035055396),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000915062237, - 0.001038062763),
    to_complex(0.004158267516, 0.003654232484),
    to_complex(- 0.000912053707, 0.001041071293),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000909043958, - 0.001044081042),
    to_complex(0.004182345566, 0.003630154434),
    to_complex(- 0.000906032932, 0.001047092068),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000903020572, - 0.001050104428),
    to_complex(0.004206444509, 0.003606055491),
    to_complex(- 0.000900006819, 0.001053118181),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000896991616, - 0.001056133384),
    to_complex(0.004230566191, 0.003581933809),
    to_complex(- 0.000893974905, 0.001059150095),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000890956628, - 0.001062168372),
    to_complex(0.004254712463, 0.003557787537),
    to_complex(- 0.000887936727, 0.001065188273),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000884915145, - 0.001068209855),
    to_complex(0.004278885183, 0.003533614817),
    to_complex(- 0.000881891821, 0.001071233179),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000878866699, - 0.001074258301),
    to_complex(0.004303086218, 0.003509413782),
    to_complex(- 0.000875839720, 0.001077285280),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000872810824, - 0.001080314176),
    to_complex(0.004327317444, 0.003485182556),
    to_complex(- 0.000869779953, 0.001083345047),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000866747048, - 0.001086377952),
    to_complex(0.004351580745, 0.003460919255),
    to_complex(- 0.000863712049, 0.001089412951),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000860674898, - 0.001092450102),
    to_complex(0.004375878016, 0.003436621984),
    to_complex(- 0.000857635534, 0.001095489466),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000854593898, - 0.001098531102),
    to_complex(0.004400211161, 0.003412288839),
    to_complex(- 0.000851549931, 0.001101575069),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000848503571, - 0.001104621429),
    to_complex(0.004424582097, 0.003387917903),
    to_complex(- 0.000845454760, 0.001107670240),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000842403435, - 0.001110721565),
    to_complex(0.004448992751, 0.003363507249),
    to_complex(- 0.000839349538, 0.001113775462),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000836293007, - 0.001116831993),
    to_complex(0.004473445064, 0.003339054936),
    to_complex(- 0.000833233780, 0.001119891220),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000830171797, - 0.001122953203),
    to_complex(0.004497940987, 0.003314559013),
    to_complex(- 0.000827106997, 0.001126018003),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000824039317, - 0.001129085683),
    to_complex(0.004522482487, 0.003290017513),
    to_complex(- 0.000820968696, 0.001132156304),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000817895072, - 0.001135229928),
    to_complex(0.004547071545, 0.003265428455),
    to_complex(- 0.000814818381, 0.001138306619),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000811738563, - 0.001141386437),
    to_complex(0.004571710157, 0.003240789843),
    to_complex(- 0.000808655553, 0.001144469447),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000805569289, - 0.001147555711),
    to_complex(0.004596400332, 0.003216099668),
    to_complex(- 0.000802479708, 0.001150645292),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000799386745, - 0.001153738255),
    to_complex(0.004621144099, 0.003191355901),
    to_complex(- 0.000796290337, 0.001156834663),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000793190419, - 0.001159934581),
    to_complex(0.004645943501, 0.003166556499),
    to_complex(- 0.000790086929, 0.001163038071),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000786979799, - 0.001166145201),
    to_complex(0.004670800600, 0.003141699400),
    to_complex(- 0.000783868967, 0.001169256033),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000780754365, - 0.001172370635),
    to_complex(0.004695717476, 0.003116782524),
    to_complex(- 0.000777635930, 0.001175489070),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000774513594, - 0.001178611406),
    to_complex(0.004720696228, 0.003091803772),
    to_complex(- 0.000771387292, 0.001181737708),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000768256957, - 0.001184868043),
    to_complex(0.004745738975, 0.003066761025),
    to_complex(- 0.000765122522, 0.001188002478),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000761983921, - 0.001191141079),
    to_complex(0.004770847856, 0.003041652144),
    to_complex(- 0.000758841084, 0.001194283916),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000755693946, - 0.001197431054),
    to_complex(0.004796025031, 0.003016474969),
    to_complex(- 0.000752542437, 0.001200582563),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000749386489, - 0.001203738511),
    to_complex(0.004821272684, 0.002991227316),
    to_complex(- 0.000746226033, 0.001206898967),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000743061000, - 0.001210064000),
    to_complex(0.004846593020, 0.002965906980),
    to_complex(- 0.000739891320, 0.001213233680),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000736716922, - 0.001216408078),
    to_complex(0.004871988269, 0.002940511731),
    to_complex(- 0.000733537738, 0.001219587262),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000730353695, - 0.001222771305),
    to_complex(0.004897460683, 0.002915039317),
    to_complex(- 0.000727164722, 0.001225960278),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000723970749, - 0.001229154251),
    to_complex(0.004923012543, 0.002889487457),
    to_complex(- 0.000720771702, 0.001232353298),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000717567510, - 0.001235557490),
    to_complex(0.004948646153, 0.002863853847),
    to_complex(- 0.000714358099, 0.001238766901),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000711143397, - 0.001241981603),
    to_complex(0.004974363847, 0.002838136153),
    to_complex(- 0.000707923329, 0.001245201671),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000704697821, - 0.001248427179),
    to_complex(0.005000167984, 0.002812332016),
    to_complex(- 0.000701466799, 0.001251658201),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000698230187, - 0.001254894813),
    to_complex(0.005026060955, 0.002786439045),
    to_complex(- 0.000694987910, 0.001258137090),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000691739891, - 0.001261385109),
    to_complex(0.005052045179, 0.002760454821),
    to_complex(- 0.000688486055, 0.001264638945),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000685226324, - 0.001267898676),
    to_complex(0.005078123106, 0.002734376894),
    to_complex(- 0.000681960620, 0.001271164380),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000678688866, - 0.001274436134),
    to_complex(0.005104297219, 0.002708202781),
    to_complex(- 0.000675410983, 0.001277714017),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000672126891, - 0.001280998109),
    to_complex(0.005130570032, 0.002681929968),
    to_complex(- 0.000668836511, 0.001284288489),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000665539764, - 0.001287585236),
    to_complex(0.005156944094, 0.002655555906),
    to_complex(- 0.000662236567, 0.001290888433),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000658926840, - 0.001294198160),
    to_complex(0.005183421990, 0.002629078010),
    to_complex(- 0.000655610501, 0.001297514499),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000652287468, - 0.001300837532),
    to_complex(0.005210006339, 0.002602493661),
    to_complex(- 0.000648957657, 0.001304167343),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000645620985, - 0.001307504015),
    to_complex(0.005236699800, 0.002575800200),
    to_complex(- 0.000642277368, 0.001310847632),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000638926720, - 0.001314198280),
    to_complex(0.005263505067, 0.002548994933),
    to_complex(- 0.000635568957, 0.001317556043),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000632203992, - 0.001320921008),
    to_complex(0.005290424876, 0.002522075124),
    to_complex(- 0.000628831738, 0.001324293262),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000625452108, - 0.001327672892),
    to_complex(0.005317462002, 0.002495037998),
    to_complex(- 0.000622065014, 0.001331059986),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000618670367, - 0.001334454633),
    to_complex(0.005344619264, 0.002467880736),
    to_complex(- 0.000615268079, 0.001337856921),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000611858058, - 0.001341266942),
    to_complex(0.005371899523, 0.002440600477),
    to_complex(- 0.000608440214, 0.001344684786),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000605014455, - 0.001348110545),
    to_complex(0.005399305685, 0.002413194315),
    to_complex(- 0.000601580689, 0.001351544311),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000598138824, - 0.001354986176),
    to_complex(0.005426840701, 0.002385659299),
    to_complex(- 0.000594688765, 0.001358436235),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000591230419, - 0.001361894581),
    to_complex(0.005454507570, 0.002357992430),
    to_complex(- 0.000587763689, 0.001365361311),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000584288479, - 0.001368836521),
    to_complex(0.005482309341, 0.002330190659),
    to_complex(- 0.000580804694, 0.001372320306),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000577312235, - 0.001375812765),
    to_complex(0.005510249111, 0.002302250889),
    to_complex(- 0.000573811004, 0.001379313996),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000570300902, - 0.001382824098),
    to_complex(0.005538330030, 0.002274169970),
    to_complex(- 0.000566781828, 0.001386343172),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000563253682, - 0.001389871318),
    to_complex(0.005566555301, 0.002245944699),
    to_complex(- 0.000559716361, 0.001393408639),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000556169764, - 0.001396955236),
    to_complex(0.005594928182, 0.002217571818),
    to_complex(- 0.000552613787, 0.001400511213),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000549048324, - 0.001404076676),
    to_complex(0.005623451988, 0.002189048012),
    to_complex(- 0.000545473271, 0.001407651729),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000541888522, - 0.001411236478),
    to_complex(0.005652130090, 0.002160369910),
    to_complex(- 0.000538293969, 0.001414831031),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000534689503, - 0.001418435497),
    to_complex(0.005680965922, 0.002131534078),
    to_complex(- 0.000531075017, 0.001422049983),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000527450399, - 0.001425674601),
    to_complex(0.005709962977, 0.002102537023),
    to_complex(- 0.000523815538, 0.001429309462),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000520170323, - 0.001432954677),
    to_complex(0.005739124814, 0.002073375186),
    to_complex(- 0.000516514639, 0.001436610361),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000512848373, - 0.001440276627),
    to_complex(0.005768455057, 0.002044044943),
    to_complex(- 0.000509171410, 0.001443953590),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000505483632, - 0.001447641368),
    to_complex(0.005797957395, 0.002014542605),
    to_complex(- 0.000501784923, 0.001451340077),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000498075163, - 0.001455049837),
    to_complex(0.005827635590, 0.001984864410),
    to_complex(- 0.000494354234, 0.001458770766),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000490622014, - 0.001462502986),
    to_complex(0.005857493473, 0.001955006527),
    to_complex(- 0.000486878381, 0.001466246619),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000483123212, - 0.001470001788),
    to_complex(0.005887534950, 0.001924965050),
    to_complex(- 0.000479356382, 0.001473768618),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000475577767, - 0.001477547233),
    to_complex(0.005917764003, 0.001894735997),
    to_complex(- 0.000471787238, 0.001481337762),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000467984668, - 0.001485140332),
    to_complex(0.005948184692, 0.001864315308),
    to_complex(- 0.000464169927, 0.001488955073),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000460342885, - 0.001492782115),
    to_complex(0.005978801159, 0.001833698841),
    to_complex(- 0.000456503410, 0.001496621590),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000452651369, - 0.001500473631),
    to_complex(0.006009617626, 0.001802882374),
    to_complex(- 0.000448786626, 0.001504338374),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000444909046, - 0.001508215954),
    to_complex(0.006040638403, 0.001771861597),
    to_complex(- 0.000441018491, 0.001512106509),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000437114823, - 0.001516010177),
    to_complex(0.006071867889, 0.001740632111),
    to_complex(- 0.000433197901, 0.001519927099),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000429267584, - 0.001523857416),
    to_complex(0.006103310573, 0.001709189427),
    to_complex(- 0.000425323727, 0.001527801273),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000421366188, - 0.001531758812),
    to_complex(0.006134971036, 0.001677528964),
    to_complex(- 0.000417394818, 0.001535730182),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000413409472, - 0.001539715528),
    to_complex(0.006166853960, 0.001645646040),
    to_complex(- 0.000409409998, 0.001543715002),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000405396247, - 0.001547728753),
    to_complex(0.006198964122, 0.001613535878),
    to_complex(- 0.000401368065, 0.001551756935),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000397325299, - 0.001555799701),
    to_complex(0.006231306405, 0.001581193595),
    to_complex(- 0.000393267793, 0.001559857207),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000389195389, - 0.001563929611),
    to_complex(0.006263885798, 0.001548614202),
    to_complex(- 0.000385107928, 0.001568017072),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000381005248, - 0.001572119752),
    to_complex(0.006296707398, 0.001515792602),
    to_complex(- 0.000376887187, 0.001576237813),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000372753581, - 0.001580371419),
    to_complex(0.006329776414, 0.001482723586),
    to_complex(- 0.000368604263, 0.001584520737),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000364439064, - 0.001588685936),
    to_complex(0.006363098175, 0.001449401825),
    to_complex(- 0.000360257814, 0.001592867186),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000356060342, - 0.001597064658),
    to_complex(0.006396678127, 0.001415821873),
    to_complex(- 0.000351846473, 0.001601278527),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000347616031, - 0.001605508969),
    to_complex(0.006430521840, 0.001381978160),
    to_complex(- 0.000343368838, 0.001609756162),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000339104715, - 0.001614020285),
    to_complex(0.006464635014, 0.001347864986),
    to_complex(- 0.000334823477, 0.001618301523),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000330524943, - 0.001622600057),
    to_complex(0.006499023479, 0.001313476521),
    to_complex(- 0.000326208924, 0.001626916076),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000321875232, - 0.001631249768),
    to_complex(0.006533693201, 0.001278806799),
    to_complex(- 0.000317523677, 0.001635601323),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000313154065, - 0.001639970935),
    to_complex(0.006568650290, 0.001243849710),
    to_complex(- 0.000308766202, 0.001644358798),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000304359888, - 0.001648765112),
    to_complex(0.006603900998, 0.001208599002),
    to_complex(- 0.000299934925, 0.001653190075),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000295491109, - 0.001657633891),
    to_complex(0.006639451728, 0.001173048272),
    to_complex(- 0.000291028237, 0.001662096763),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000286546099, - 0.001666578901),
    to_complex(0.006675309038, 0.001137190962),
    to_complex(- 0.000282044487, 0.001671080513),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000277523188, - 0.001675601812),
    to_complex(0.006711479646, 0.001101020354),
    to_complex(- 0.000272981986, 0.001680143014),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000268420665, - 0.001684704335),
    to_complex(0.006747970437, 0.001064529563),
    to_complex(- 0.000263839003, 0.001689285997),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000259236778, - 0.001693888222),
    to_complex(0.006784788465, 0.001027711535),
    to_complex(- 0.000254613763, 0.001698511237),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000249969730, - 0.001703155270),
    to_complex(0.006821940963, 0.000990559037),
    to_complex(- 0.000245304447, 0.001707820553),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000240617679, - 0.001712507321),
    to_complex(0.006859435344, 0.000953064656),
    to_complex(- 0.000235909189, 0.001717215811),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000231178736, - 0.001721946264),
    to_complex(0.006897279213, 0.000915220787),
    to_complex(- 0.000226426076, 0.001726698924),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000221650963, - 0.001731474037),
    to_complex(0.006935480368, 0.000877019632),
    to_complex(- 0.000216853146, 0.001736271854),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000212032373, - 0.001741092627),
    to_complex(0.006974046811, 0.000838453189),
    to_complex(- 0.000207188386, 0.001745936614),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000202320926, - 0.001750804074),
    to_complex(0.007012986754, 0.000799513246),
    to_complex(- 0.000197429730, 0.001755695270),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000192514530, - 0.001760610470),
    to_complex(0.007052308623, 0.000760191377),
    to_complex(- 0.000187575056, 0.001765549944),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000182611035, - 0.001770513965),
    to_complex(0.007092021070, 0.000720478930),
    to_complex(- 0.000177622189, 0.001775502811),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000172608236, - 0.001780516764),
    to_complex(0.007132132978, 0.000680367022),
    to_complex(- 0.000167568891, 0.001785556109),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000162503866, - 0.001790621134),
    to_complex(0.007172653473, 0.000639846527),
    to_complex(- 0.000157412867, 0.001795712133),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000152295598, - 0.001800829402),
    to_complex(0.007213591927, 0.000598908073),
    to_complex(- 0.000147151758, 0.001805973242),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000141981041, - 0.001811143959),
    to_complex(0.007254957972, 0.000557542028),
    to_complex(- 0.000136783138, 0.001816341862),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000131557736, - 0.001821567264),
    to_complex(0.007296761505, 0.000515738495),
    to_complex(- 0.000126304517, 0.001826820483),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000121023158, - 0.001832101842),
    to_complex(0.007339012703, 0.000473487297),
    to_complex(- 0.000115713333, 0.001837411667),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000110374709, - 0.001842750291),
    to_complex(0.007381722029, 0.000430777971),
    to_complex(- 0.000105006951, 0.001848118049),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000099609717, - 0.001853515283),
    to_complex(0.007424900242, 0.000387599758),
    to_complex(- 0.000094182663, 0.001858942337),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000088725436, - 0.001864399564),
    to_complex(0.007468558414, 0.000343941586),
    to_complex(- 0.000083237681, 0.001869887319),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000077719036, - 0.001875405964),
    to_complex(0.007512707934, 0.000299792066),
    to_complex(- 0.000072169137, 0.001880955863),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000066587610, - 0.001886537390),
    to_complex(0.007557360525, 0.000255139475),
    to_complex(- 0.000060974079, 0.001892150921),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000055328161, - 0.001897796839),
    to_complex(0.007602528255, 0.000209971745),
    to_complex(- 0.000049649468, 0.001903475532),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000043937606, - 0.001909187394),
    to_complex(0.007648223552, 0.000164276448),
    to_complex(- 0.000038192175, 0.001914932825),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000032412769, - 0.001920712231),
    to_complex(0.007694459215, 0.000118040785),
    to_complex(- 0.000026598975, 0.001926526025),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000020750376, - 0.001932374624),
    to_complex(0.007741248430, 0.000071251570),
    to_complex(- 0.000014866548, 0.001938258452),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000008947058, - 0.001944177942),
    to_complex(0.007788604785, 0.000023895215),
    to_complex(- 0.000002991470, 0.001950133530),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.000003000662, - 0.001956125662),
    to_complex(0.007836542286, - 0.000024042286),
    to_complex(0.000009029787, 0.001962154787),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.000015096365, - 0.001968221365),
    to_complex(0.007885075374, - 0.000072575374),
    to_complex(0.000021200860, 0.001974325860),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.000027343746, - 0.001980468746),
    to_complex(0.007934218942, - 0.000121718942),
    to_complex(0.000033525503, 0.001986650503),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.000039746617, - 0.001992871617),
    to_complex(0.007983988351, - 0.000171488351),
    to_complex(0.000046007584, 0.001999132584),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.000052308908, - 0.002005433908),
    to_complex(0.008034399454, - 0.000221899454),
    to_complex(0.000058651100, 0.002011776100),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.000065034679, - 0.002018159679),
    to_complex(0.008085468613, - 0.000272968613),
    to_complex(0.000071460173, 0.002024585173),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.000077928118, - 0.002031053118),
    to_complex(0.008137212718, - 0.000324712718),
    to_complex(0.000084439059, 0.002037564059),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.000090993551, - 0.002044118551),
    to_complex(0.008189649215, - 0.000377149215),
    to_complex(0.000097592156, 0.002050717156),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.000104235447, - 0.002057360447),
    to_complex(0.008242796122, - 0.000430296122),
    to_complex(0.000110924005, 0.002064049005),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.000117658422, - 0.002070783422),
    to_complex(0.008296672060, - 0.000484172060),
    to_complex(0.000124439299, 0.002077564299),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.000131267248, - 0.002084392248),
    to_complex(0.008351296274, - 0.000538796274),
    to_complex(0.000138142891, 0.002091267891),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.000145066859, - 0.002098191859),
    to_complex(0.008406688662, - 0.000594188662),
    to_complex(0.000152039796, 0.002105164796),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.000159062355, - 0.002112187355),
    to_complex(0.008462869804, - 0.000650369804),
    to_complex(0.000166135203, 0.002119260203),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.000173259015, - 0.002126384015),
    to_complex(0.008519860990, - 0.000707360990),
    to_complex(0.000180434480, 0.002133559480),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.000187662299, - 0.002140787299),
    to_complex(0.008577684251, - 0.000765184251),
    to_complex(0.000194943183, 0.002148068183),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.000202277859, - 0.002155402859),
    to_complex(0.008636362396, - 0.000823862396),
    to_complex(0.000209667064, 0.002162792064),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.000217111549, - 0.002170236549),
    to_complex(0.008695919041, - 0.000883419041),
    to_complex(0.000224612079, 0.002177737079),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.000232169431, - 0.002185294431),
    to_complex(0.008756378651, - 0.000943878651),
    to_complex(0.000239784398, 0.002192909398),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.000247457786, - 0.002200582786),
    to_complex(0.008817766576, - 0.001005266576),
    to_complex(0.000255190416, 0.002208315416),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.000262983124, - 0.002216108124),
    to_complex(0.008880109092, - 0.001067609092),
    to_complex(0.000270836762, 0.002223961762),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.000278752196, - 0.002231877196),
    to_complex(0.008943433446, - 0.001130933446),
    to_complex(0.000286730309, 0.002239855309),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.000294772001, - 0.002247897001),
    to_complex(0.009007767898, - 0.001195267898),
    to_complex(0.000302878188, 0.002256003188),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.000311049804, - 0.002264174804),
    to_complex(0.009073141774, - 0.001260641774),
    to_complex(0.000319287799, 0.002272412799),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.000327593143, - 0.002280718143),
    to_complex(0.009139585514, - 0.001327085514),
    to_complex(0.000335966823, 0.002289091823),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.000344409846, - 0.002297534846),
    to_complex(0.009207130723, - 0.001394630723),
    to_complex(0.000352923238, 0.002306048238),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.000361508044, - 0.002314633044),
    to_complex(0.009275810237, - 0.001463310237),
    to_complex(0.000370165330, 0.002323290330),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.000378896183, - 0.002332021183),
    to_complex(0.009345658172, - 0.001533158172),
    to_complex(0.000387701712, 0.002340826712),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.000396583046, - 0.002349708046),
    to_complex(0.009416709999, - 0.001604209999),
    to_complex(0.000405541339, 0.002358666339),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.000414577764, - 0.002367702764),
    to_complex(0.009489002604, - 0.001676502604),
    to_complex(0.000423693523, 0.002376818523),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.000432889836, - 0.002386014836),
    to_complex(0.009562574363, - 0.001750074363),
    to_complex(0.000442167954, 0.002395292954),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.000451529149, - 0.002404654149),
    to_complex(0.009637465219, - 0.001824965219),
    to_complex(0.000460974720, 0.002414099720),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.000470505993, - 0.002423630993),
    to_complex(0.009713716762, - 0.001901216762),
    to_complex(0.000480124323, 0.002433249323),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.000489831091, - 0.002442956091),
    to_complex(0.009791372317, - 0.001978872317),
    to_complex(0.000499627708, 0.002452752708),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.000509515614, - 0.002462640614),
    to_complex(0.009870477034, - 0.002057977034),
    to_complex(0.000519496279, 0.002472621279),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.000529571207, - 0.002482696207),
    to_complex(0.009951077986, - 0.002138577986),
    to_complex(0.000539741930, 0.002492866930),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.000550010015, - 0.002503135015),
    to_complex(0.010033224273, - 0.002220724273),
    to_complex(0.000560377065, 0.002513502065),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.000570844714, - 0.002523969714),
    to_complex(0.010116967136, - 0.002304467136),
    to_complex(0.000581414634, 0.002534539634),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.000592088532, - 0.002545213532),
    to_complex(0.010202360070, - 0.002389860070),
    to_complex(0.000602868155, 0.002555993155),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.000613755288, - 0.002566880288),
    to_complex(0.010289458953, - 0.002476958953),
    to_complex(0.000624751754, 0.002577876754),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.000635859419, - 0.002588984419),
    to_complex(0.010378322181, - 0.002565822181),
    to_complex(0.000647080190, 0.002600205190),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.000658416020, - 0.002611541020),
    to_complex(0.010469010811, - 0.002656510811),
    to_complex(0.000669868902, 0.002622993902),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.000681440879, - 0.002634565879),
    to_complex(0.010561588717, - 0.002749088717),
    to_complex(0.000693134040, 0.002646259040),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.000704950520, - 0.002658075520),
    to_complex(0.010656122748, - 0.002843622748),
    to_complex(0.000716892508, 0.002670017508),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.000728962243, - 0.002682087243),
    to_complex(0.010752682915, - 0.002940182915),
    to_complex(0.000741162015, 0.002694287015),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.000753494172, - 0.002706619172),
    to_complex(0.010851342571, - 0.003038842571),
    to_complex(0.000765961115, 0.002719086115),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.000778565306, - 0.002731690306),
    to_complex(0.010952178618, - 0.003139678618),
    to_complex(0.000791309265, 0.002744434265),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.000804195572, - 0.002757320572),
    to_complex(0.011055271724, - 0.003242771724),
    to_complex(0.000817226874, 0.002770351874),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.000830405881, - 0.002783530881),
    to_complex(0.011160706556, - 0.003348206556),
    to_complex(0.000843735370, 0.002796860370),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.000857218190, - 0.002810343190),
    to_complex(0.011268572034, - 0.003456072034),
    to_complex(0.000870857260, 0.002823982260),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.000884655572, - 0.002837780572),
    to_complex(0.011378961600, - 0.003566461600),
    to_complex(0.000898616196, 0.002851741196),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.000912742281, - 0.002865867281),
    to_complex(0.011491973509, - 0.003679473509),
    to_complex(0.000927037056, 0.002880162056),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.000941503836, - 0.002894628836),
    to_complex(0.011607711147, - 0.003795211147),
    to_complex(0.000956146021, 0.002909271021),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.000970967100, - 0.002924092100),
    to_complex(0.011726283367, - 0.003913783367),
    to_complex(0.000985970658, 0.002939095658),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.001001160372, - 0.002954285372),
    to_complex(0.011847804858, - 0.004035304858),
    to_complex(0.001016540021, 0.002969665021),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.001032113483, - 0.002985238483),
    to_complex(0.011972396542, - 0.004159896542),
    to_complex(0.001047884745, 0.003001009745),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.001063857902, - 0.003016982902),
    to_complex(0.012100186005, - 0.004287686005),
    to_complex(0.001080037162, 0.003033162162),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.001096426850, - 0.003049551850),
    to_complex(0.012231307960, - 0.004418807960),
    to_complex(0.001113031414, 0.003066156414),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.001129855426, - 0.003082980426),
    to_complex(0.012365904754, - 0.004553404754),
    to_complex(0.001146903587, 0.003100028587),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.001164180736, - 0.003117305736),
    to_complex(0.012504126920, - 0.004691626920),
    to_complex(0.001181691848, 0.003134816848),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.001199442046, - 0.003152567046),
    to_complex(0.012646133770, - 0.004833633770),
    to_complex(0.001217436599, 0.003170561599),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.001235680936, - 0.003188805936),
    to_complex(0.012792094048, - 0.004979594048),
    to_complex(0.001254180643, 0.003207305643),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.001272941476, - 0.003226066476),
    to_complex(0.012942186641, - 0.005129686641),
    to_complex(0.001291969363, 0.003245094363),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.001311270415, - 0.003264395415),
    to_complex(0.013096601347, - 0.005284101347),
    to_complex(0.001330850926, 0.003283975926),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.001350717387, - 0.003303842387),
    to_complex(0.013255539729, - 0.005443039729),
    to_complex(0.001370876491, 0.003324001491),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.001391335139, - 0.003344460139),
    to_complex(0.013419216035, - 0.005606716035),
    to_complex(0.001412100452, 0.003365225452),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.001433179777, - 0.003386304777),
    to_complex(0.013587858215, - 0.005775358215),
    to_complex(0.001454580696, 0.003407705696),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.001476311039, - 0.003429436039),
    to_complex(0.013761709038, - 0.005949209038),
    to_complex(0.001498378888, 0.003451503888),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.001520792594, - 0.003473917594),
    to_complex(0.013941027311, - 0.006128527311),
    to_complex(0.001543560783, 0.003496685783),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.001566692372, - 0.003519817372),
    to_complex(0.014126089233, - 0.006313589233),
    to_complex(0.001590196575, 0.003543321575),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.001614082923, - 0.003567207923),
    to_complex(0.014317189876, - 0.006504689876),
    to_complex(0.001638361273, 0.003591486273),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.001663041823, - 0.003616166823),
    to_complex(0.014514644829, - 0.006702144829),
    to_complex(0.001688135127, 0.003641260127),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.001713652112, - 0.003666777112),
    to_complex(0.014718792015, - 0.006906292015),
    to_complex(0.001739604090, 0.003692729090),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.001766002783, - 0.003719127783),
    to_complex(0.014929993699, - 0.007117493699),
    to_complex(0.001792860334, 0.003745985334),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.001820189331, - 0.003773314331),
    to_complex(0.015148638727, - 0.007336138727),
    to_complex(0.001848002826, 0.003801127826),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.001876314355, - 0.003829439355),
    to_complex(0.015375145004, - 0.007562645004),
    to_complex(0.001905137964, 0.003858262964),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.001934488230, - 0.003887613230),
    to_complex(0.015609962267, - 0.007797462267),
    to_complex(0.001964380289, 0.003917505289),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.001994829860, - 0.003947954860),
    to_complex(0.015853575171, - 0.008041075171),
    to_complex(0.002025853278, 0.003978978278),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.002057467519, - 0.004010592519),
    to_complex(0.016106506750, - 0.008294006750),
    to_complex(0.002089690236, 0.004042815236),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.002122539791, - 0.004075664791),
    to_complex(0.016369322293, - 0.008556822293),
    to_complex(0.002156035291, 0.004109160291),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.002190196627, - 0.004143321627),
    to_complex(0.016642633696, - 0.008830133696),
    to_complex(0.002225044515, 0.004178169515),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.002260600538, - 0.004213725538),
    to_complex(0.016927104375, - 0.009114604375),
    to_complex(0.002296887193, 0.004250012193),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.002333927938, - 0.004287052938),
    to_complex(0.017223454802, - 0.009410954802),
    to_complex(0.002371747245, 0.004324872245),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.002410370658, - 0.004363495658),
    to_complex(0.017532468773, - 0.009719968773),
    to_complex(0.002449824848, 0.004402949848),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.002490137678, - 0.004443262678),
    to_complex(0.017855000528, - 0.010042500528),
    to_complex(0.002531338269, 0.004484463269),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.002573457077, - 0.004526582077),
    to_complex(0.018191982843, - 0.010379482843),
    to_complex(0.002616525961, 0.004569650961),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.002660578275, - 0.004613703275),
    to_complex(0.018544436275, - 0.010731936275),
    to_complex(0.002705648947, 0.004658773947),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.002751774583, - 0.004704899583),
    to_complex(0.018913479732, - 0.011100979732),
    to_complex(0.002798993560, 0.004752118560),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.002847346139, - 0.004800471139),
    to_complex(0.019300342622, - 0.011487842622),
    to_complex(0.002896874583, 0.004849999583),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.002947623279, - 0.004900748279),
    to_complex(0.019706378832, - 0.011893878832),
    to_complex(0.002999638878, 0.004952763878),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.003052970435, - 0.005006095435),
    to_complex(0.020133082903, - 0.012320582903),
    to_complex(0.003107669574, 0.005060794574),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.003163790650, - 0.005116915650),
    to_complex(0.020582108778, - 0.012769608778),
    to_complex(0.003221390940, 0.005174515940),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.003280530834, - 0.005233655834),
    to_complex(0.021055291641, - 0.013242791641),
    to_complex(0.003341274056, 0.005294399056),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.003403687895, - 0.005356812895),
    to_complex(0.021554673440, - 0.013742173440),
    to_complex(0.003467843456, 0.005420968456),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.003533815938, - 0.005486940938),
    to_complex(0.022082532858, - 0.014270032858),
    to_complex(0.003601684928, 0.005554809928),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.003671534732, - 0.005624659732),
    to_complex(0.022641420645, - 0.014828920645),
    to_complex(0.003743454726, 0.005696579726),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.003817539744, - 0.005770664744),
    to_complex(0.023234201470, - 0.015421701470),
    to_complex(0.003893890499, 0.005847015499),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.003972614051, - 0.005925739051),
    to_complex(0.023864103757, - 0.016051603757),
    to_complex(0.004053824308, 0.006006949308),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.004137642590, - 0.006090767590),
    to_complex(0.024534779311, - 0.016722279311),
    to_complex(0.004224198236, 0.006177323236),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.004313629280, - 0.006266754280),
    to_complex(0.025250375081, - 0.017437875081),
    to_complex(0.004406083193, 0.006359208193),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.004501717707, - 0.006454842707),
    to_complex(0.026015620025, - 0.018203120025),
    to_complex(0.004600701718, 0.006553826718),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.004703216296, - 0.006656341296),
    to_complex(0.026835930933, - 0.019023430933),
    to_complex(0.004809455801, 0.006762580801),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.004919629121, - 0.006872754121),
    to_complex(0.027717542202, - 0.019905042202),
    to_complex(0.005033961062, 0.006987086062),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.005152693889, - 0.007105818889),
    to_complex(0.028667666156, - 0.020855166156),
    to_complex(0.005276089058, 0.007229214058),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.005404429149, - 0.007357554149),
    to_complex(0.029694692621, - 0.021882192621),
    to_complex(0.005538020051, 0.007491145051),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.005677193408, - 0.007630318408),
    to_complex(0.030808439456, - 0.022995939456),
    to_complex(0.005822309394, 0.007775434394),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.005973759849, - 0.007926884849),
    to_complex(0.032020469896, - 0.024207969896),
    to_complex(0.006131971829, 0.008085096829),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.006297411662, - 0.008250536662),
    to_complex(0.033344498452, - 0.025531998452),
    to_complex(0.006470589566, 0.008423714566),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.006652064936, - 0.008605189936),
    to_complex(0.034796915612, - 0.026984415612),
    to_complex(0.006842452413, 0.008795577413),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.007042428882, - 0.008995553882),
    to_complex(0.036397473994, - 0.028584973994),
    to_complex(0.007252741554, 0.009205866554),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.007474217340, - 0.009427342340),
    to_complex(0.038170197021, - 0.030357697021),
    to_complex(0.007707773773, 0.009660898773),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.007954431767, - 0.009907556767),
    to_complex(0.040144599158, - 0.032332099158),
    to_complex(0.008215330605, 0.010168455605),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.008491745603, - 0.010444870603),
    to_complex(0.042357349863, - 0.034544849863),
    to_complex(0.008785109036, 0.010738234036),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.009097035057, - 0.011050160057),
    to_complex(0.044854581647, - 0.037042081647),
    to_complex(0.009429349511, 0.011382474511),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.009784125813, - 0.011737250813),
    to_complex(0.047695153199, - 0.039882653199),
    to_complex(0.010163728385, 0.012116853385),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.010570865562, - 0.012523990562),
    to_complex(0.050955362780, - 0.043142862780),
    to_complex(0.011008654486, 0.012961779486),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.011480701260, - 0.013433826260),
    to_complex(0.054735924060, - 0.046923424060),
    to_complex(0.011991200739, 0.013944325739),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.012545061796, - 0.014498186796),
    to_complex(0.059172581505, - 0.051360081505),
    to_complex(0.013148065990, 0.015101190990),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.013807070518, - 0.015760195518),
    to_complex(0.064452791713, - 0.056640291713),
    to_complex(0.014530270569, 0.016483395569),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.015327542393, - 0.017280667393),
    to_complex(0.070842940328, - 0.063030440328),
    to_complex(0.016210897645, 0.018164022645),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.017195093499, - 0.019148218499),
    to_complex(0.078734770882, - 0.070922270882),
    to_complex(0.018298464629, 0.020251589629),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.019544077231, - 0.021497202231),
    to_complex(0.088728956729, - 0.080916456729),
    to_complex(0.020961360594, 0.022914485594),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.022588463793, - 0.024541588793),
    to_complex(0.101795816292, - 0.093983316292),
    to_complex(0.024475743603, 0.026428868603),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.026691072202, - 0.028644197202),
    to_complex(0.119611354027, - 0.111798854027),
    to_complex(0.029328177833, 0.031281302833),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.032520253260, - 0.034473378260),
    to_complex(0.145341356024, - 0.137528856024),
    to_complex(0.036463170193, 0.038416295193),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.041457265253, - 0.043410390253),
    to_complex(0.185769649482, - 0.177957149482),
    to_complex(0.047987697593, 0.049940822593),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.056892469387, - 0.058845594387),
    to_complex(0.258534184926, - 0.250721684926),
    to_complex(0.069754473622, 0.071707598622),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.089965623841, - 0.091918748841),
    to_complex(0.428307447286, - 0.420494947286),
    to_complex(0.126344895250, 0.128298020250),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.211228530259, - 0.213181655259),
    to_complex(1.277141799991, - 1.269329299991),
    to_complex(0.635642710525, 0.637595835525));

  constant INPUT_DATA_2048_16QAM_NOISY : complex_array(0 to 2047) := (-- Symbol Error Rate: 0.0019531
    to_complex(0.010090149999, 0.008979943628),
    to_complex(0.640239971539, 0.638276107866),
    to_complex(- 1.271339647715, 1.287695766422),
    to_complex(- 0.209796926272, - 0.203272630023),
    to_complex(0.000359448285, - 0.000267899362),
    to_complex(0.131210783057, 0.113188541497),
    to_complex(- 0.417978885796, 0.428821697587),
    to_complex(- 0.090098887345, - 0.092313033811),
    to_complex(- 0.007518355636, 0.002861134585),
    to_complex(0.075402087285, 0.081176366467),
    to_complex(- 0.252255006455, 0.284116375575),
    to_complex(- 0.066312905613, - 0.040697187530),
    to_complex(0.008210282822, 0.009883150262),
    to_complex(0.063979016711, 0.042725625778),
    to_complex(- 0.168711664993, 0.176920497115),
    to_complex(- 0.040081053687, - 0.048188759204),
    to_complex(- 0.002233027675, 0.003750963552),
    to_complex(0.040138077391, 0.031897895999),
    to_complex(- 0.137004714366, 0.155465729987),
    to_complex(- 0.031398552267, - 0.037111566951),
    to_complex(- 0.001819329257, 0.004779767935),
    to_complex(0.024585089881, 0.025170728226),
    to_complex(- 0.109879655483, 0.122641309839),
    to_complex(- 0.034665137760, - 0.023504408058),
    to_complex(- 0.003323710863, - 0.003133716480),
    to_complex(0.033914909882, 0.016129005229),
    to_complex(- 0.097832970576, 0.095864706012),
    to_complex(- 0.022384065099, - 0.014243127088),
    to_complex(- 0.001662116836, 0.002387013141),
    to_complex(0.018084271753, 0.015001822512),
    to_complex(- 0.080830865649, 0.095576845636),
    to_complex(- 0.022542861211, - 0.026367141428),
    to_complex(- 0.005006663411, - 0.004567012960),
    to_complex(0.016020720347, 0.021881582156),
    to_complex(- 0.060861931177, 0.067198796948),
    to_complex(- 0.014357700288, - 0.024828911342),
    to_complex(0.004668344058, - 0.000914004526),
    to_complex(0.015460518731, 0.019603626804),
    to_complex(- 0.064860708331, 0.063175745339),
    to_complex(- 0.028908403301, - 0.027862650916),
    to_complex(0.003165693949, 0.001636483649),
    to_complex(0.008687386607, 0.013294623942),
    to_complex(- 0.048735489446, 0.059585006328),
    to_complex(- 0.014529005836, - 0.011011840907),
    to_complex(- 0.001348554512, 0.001172678188),
    to_complex(0.014983803942, 0.019607349905),
    to_complex(- 0.049498361914, 0.057330976860),
    to_complex(- 0.020266610776, - 0.026719447596),
    to_complex(- 0.003226043558, 0.011893359476),
    to_complex(0.020729412875, 0.000587965459),
    to_complex(- 0.062346400473, 0.054608456715),
    to_complex(- 0.007366605134, - 0.013451584576),
    to_complex(0.007458760263, 0.003342652156),
    to_complex(0.016178480118, 0.007682900438),
    to_complex(- 0.037902367798, 0.047245268462),
    to_complex(- 0.009335918343, - 0.008628084906),
    to_complex(0.007114574487, 0.012981938868),
    to_complex(0.011946305696, - 0.000574573578),
    to_complex(- 0.047282077311, 0.041296494403),
    to_complex(- 0.014070213703, - 0.010265456432),
    to_complex(0.007686717500, 0.009213974578),
    to_complex(0.015182580103, 0.016172749894),
    to_complex(- 0.041213436001, 0.037008724451),
    to_complex(- 0.001303587461, - 0.005048784660),
    to_complex(0.000845797082, 0.004262432888),
    to_complex(0.000179383649, 0.004545328886),
    to_complex(- 0.031472314773, 0.031323972250),
    to_complex(- 0.002054674214, 0.003226359352),
    to_complex(0.010836598990, 0.004057308858),
    to_complex(0.009374901130, 0.008518141732),
    to_complex(- 0.037924563430, 0.035936644729),
    to_complex(- 0.019585920213, - 0.012695344490),
    to_complex(0.002091336102, 0.002243728766),
    to_complex(0.013698230994, - 0.000544309325),
    to_complex(- 0.024836655245, 0.043377462198),
    to_complex(- 0.012165634997, - 0.010857173970),
    to_complex(- 0.002368741944, 0.008210601255),
    to_complex(0.005335304414, 0.009388067070),
    to_complex(- 0.027576700474, 0.024581804151),
    to_complex(- 0.012221832952, 0.004580088105),
    to_complex(0.004743216649, - 0.007922476673),
    to_complex(0.008032757116, - 0.000097760418),
    to_complex(- 0.032134821617, 0.033134264231),
    to_complex(- 0.006783153853, - 0.014079587751),
    to_complex(0.004843799772, 0.002153838575),
    to_complex(0.013528909813, - 0.003569547038),
    to_complex(- 0.014818979703, 0.039089500808),
    to_complex(- 0.001260738160, - 0.002087196561),
    to_complex(- 0.001945617279, - 0.004979392976),
    to_complex(0.009992645004, 0.012407557109),
    to_complex(- 0.020131525017, 0.042746496808),
    to_complex(- 0.016332345432, - 0.012091980129),
    to_complex(0.007007248998, 0.000185659344),
    to_complex(0.003371826554, - 0.004629868008),
    to_complex(- 0.011748418607, 0.037532383995),
    to_complex(0.004151187233, 0.007354551290),
    to_complex(- 0.002553317560, 0.013576647417),
    to_complex(- 0.001225863100, 0.009542528480),
    to_complex(- 0.026180982931, 0.026314256813),
    to_complex(- 0.010080324460, - 0.024596354340),
    to_complex(0.004741250678, - 0.001798161629),
    to_complex(0.008968658953, 0.010586826248),
    to_complex(- 0.016620461851, 0.026090207401),
    to_complex(0.003696841858, - 0.010916856330),
    to_complex(- 0.000418451500, 0.008834109032),
    to_complex(0.006301369155, - 0.001199794187),
    to_complex(- 0.023471665372, 0.018346351709),
    to_complex(- 0.011206621920, - 0.008997112892),
    to_complex(0.002774146927, 0.008796928186),
    to_complex(0.011207517282, 0.011536924858),
    to_complex(- 0.021603947552, 0.020225185169),
    to_complex(- 0.007652709509, - 0.015500460664),
    to_complex(- 0.002336012760, - 0.010513610066),
    to_complex(0.006560195148, 0.018500090210),
    to_complex(- 0.022942353882, 0.026918750641),
    to_complex(- 0.008442152156, - 0.012805419817),
    to_complex(0.007666752428, 0.006126492992),
    to_complex(- 0.012950227152, 0.008087075671),
    to_complex(- 0.020350774141, 0.016841533405),
    to_complex(- 0.017133799919, - 0.003967637240),
    to_complex(0.003758889026, - 0.003614610010),
    to_complex(0.013712056381, 0.007610709837),
    to_complex(- 0.008320569579, 0.044437376376),
    to_complex(- 0.003478116050, 0.001755067632),
    to_complex(0.006272724845, 0.006273013984),
    to_complex(0.006976423583, 0.004487624311),
    to_complex(- 0.006978995324, 0.019697859443),
    to_complex(- 0.024010175949, - 0.010530635202),
    to_complex(- 0.012775199748, - 0.013079936719),
    to_complex(0.001732500336, 0.002767953722),
    to_complex(- 0.012147528654, 0.010246165797),
    to_complex(0.001560923339, - 0.000682699203),
    to_complex(0.009631285449, 0.005929710260),
    to_complex(- 0.007278264304, - 0.001197774713),
    to_complex(- 0.006034831788, 0.020152198211),
    to_complex(0.007498108030, - 0.003081794609),
    to_complex(0.000311072451, 0.006764828689),
    to_complex(- 0.004201335662, - 0.003320496525),
    to_complex(0.007122594443, 0.023772463055),
    to_complex(- 0.011512817343, - 0.006335572134),
    to_complex(0.003988501705, - 0.016386890497),
    to_complex(0.002892744965, - 0.009544531448),
    to_complex(- 0.012798688108, 0.008595485413),
    to_complex(0.007842312128, - 0.002709479525),
    to_complex(- 0.005111673691, 0.007927017678),
    to_complex(0.013067429170, - 0.003812892210),
    to_complex(- 0.001334268791, 0.013962845929),
    to_complex(0.000164610902, - 0.000033103430),
    to_complex(0.005056360102, 0.006361145264),
    to_complex(0.013973046496, 0.000998993726),
    to_complex(- 0.015378202812, 0.022209025874),
    to_complex(- 0.006749253632, - 0.002971186628),
    to_complex(- 0.003564481967, - 0.007067843692),
    to_complex(0.012487854668, 0.001537849844),
    to_complex(- 0.006241106611, 0.019746644531),
    to_complex(0.001162367035, 0.005827209027),
    to_complex(- 0.010826288634, 0.003537903445),
    to_complex(0.000403915150, 0.001811829044),
    to_complex(- 0.017324559185, 0.012351391268),
    to_complex(- 0.016156925188, 0.000151325943),
    to_complex(- 0.001771808578, - 0.010381749023),
    to_complex(0.002869727429, - 0.010703895831),
    to_complex(- 0.006288482187, 0.024642587508),
    to_complex(0.001836628924, - 0.010107218220),
    to_complex(- 0.006675010555, 0.003746026692),
    to_complex(0.006434678946, 0.006007246907),
    to_complex(- 0.013796934767, 0.025602538479),
    to_complex(- 0.002048017627, - 0.005322085151),
    to_complex(0.009851484025, 0.004255642395),
    to_complex(- 0.004288357399, 0.005007003474),
    to_complex(- 0.010684713045, 0.034277734662),
    to_complex(- 0.000969993313, 0.003678383770),
    to_complex(- 0.011983321983, - 0.003508713856),
    to_complex(0.012370754175, - 0.001894552330),
    to_complex(- 0.008129574488, 0.019804953253),
    to_complex(0.012593038306, 0.002787862558),
    to_complex(0.005978556466, - 0.001438884824),
    to_complex(0.010087362394, - 0.002884752736),
    to_complex(0.000886828545, 0.029549774773),
    to_complex(- 0.006613011237, - 0.002637522261),
    to_complex(0.008308817766, - 0.012771343537),
    to_complex(0.003399290486, - 0.012984581997),
    to_complex(- 0.005562540769, 0.019989412678),
    to_complex(- 0.003296346426, - 0.005018357940),
    to_complex(- 0.002014225133, 0.007635091838),
    to_complex(- 0.002717886176, 0.003588953662),
    to_complex(- 0.009404391120, 0.018980074570),
    to_complex(- 0.003476904929, 0.004505822923),
    to_complex(0.000329515508, - 0.004831867077),
    to_complex(0.004436105925, 0.002857724207),
    to_complex(- 0.010638934876, 0.019586470448),
    to_complex(- 0.000132791428, 0.003141362092),
    to_complex(0.005273563514, 0.013391481614),
    to_complex(0.010163626542, 0.005445631115),
    to_complex(- 0.008983541801, 0.012006031240),
    to_complex(- 0.007753551639, - 0.003991945234),
    to_complex(0.011352784728, - 0.005220394583),
    to_complex(0.002920351923, 0.007812248228),
    to_complex(- 0.011546101414, 0.016813629606),
    to_complex(- 0.009429611180, - 0.014561836606),
    to_complex(- 0.000859419817, 0.003744240195),
    to_complex(0.004460167943, 0.005000893674),
    to_complex(- 0.011062294327, 0.026128338536),
    to_complex(- 0.004641676533, - 0.002274917546),
    to_complex(- 0.008714062132, - 0.000878977360),
    to_complex(- 0.000669593222, 0.005511639744),
    to_complex(- 0.016026351612, 0.022772828229),
    to_complex(- 0.003698362626, - 0.005770719774),
    to_complex(0.006423680888, - 0.011826695593),
    to_complex(- 0.000101544072, 0.008051779422),
    to_complex(- 0.014117785813, 0.004583489084),
    to_complex(- 0.011305337458, - 0.000962478204),
    to_complex(0.003885470346, 0.004465497595),
    to_complex(0.005526348993, 0.002783650840),
    to_complex(- 0.006563557153, 0.022950721926),
    to_complex(0.004115735886, - 0.003562983268),
    to_complex(- 0.010647709888, - 0.002567319559),
    to_complex(0.013444190923, 0.000225435333),
    to_complex(- 0.018550837349, 0.009819649027),
    to_complex(0.003547932977, 0.005808827507),
    to_complex(0.001659017860, - 0.000098302306),
    to_complex(0.000007938315, 0.004733891781),
    to_complex(- 0.002446022379, 0.015182971148),
    to_complex(0.002637183474, 0.012153235696),
    to_complex(- 0.001743830282, 0.005506534955),
    to_complex(0.009896350787, 0.001663790344),
    to_complex(0.004977208353, 0.027487227328),
    to_complex(0.004089586762, - 0.001751561664),
    to_complex(0.009891048232, 0.002667116448),
    to_complex(- 0.002525953399, - 0.000263074220),
    to_complex(- 0.014634299467, 0.015815009699),
    to_complex(- 0.016377581028, - 0.008418415108),
    to_complex(0.006861499089, 0.009758046453),
    to_complex(- 0.002054307185, 0.008163222751),
    to_complex(- 0.012734725764, 0.020123633648),
    to_complex(- 0.011880226748, 0.003230784835),
    to_complex(- 0.001574200468, 0.004476726466),
    to_complex(- 0.000102846551, 0.005417550886),
    to_complex(- 0.004745481333, 0.009588290671),
    to_complex(- 0.010945325664, - 0.007668541554),
    to_complex(- 0.002182835209, - 0.015853761720),
    to_complex(0.004554814583, 0.005772853235),
    to_complex(0.005288411966, 0.012701623248),
    to_complex(0.005168364902, - 0.004802166668),
    to_complex(- 0.002283011883, 0.004092244161),
    to_complex(0.014458539370, 0.025006586722),
    to_complex(0.001120678581, 0.001737962930),
    to_complex(- 0.009342755218, - 0.014322091999),
    to_complex(- 0.004188396652, - 0.004688890408),
    to_complex(0.001444232053, - 0.000586159408),
    to_complex(0.004342410243, 0.003650815118),
    to_complex(- 0.005299065921, - 0.015435311287),
    to_complex(0.009109006689, - 0.010765324041),
    to_complex(0.002667176951, 0.009676073036),
    to_complex(0.009071821280, 0.004984648083),
    to_complex(0.008234017400, - 0.006568854685),
    to_complex(- 0.013363866501, - 0.009375841176),
    to_complex(0.009516440378, 0.010392761530),
    to_complex(- 0.009023529186, 0.005674577115),
    to_complex(- 0.014746624593, - 0.004674627045),
    to_complex(- 0.004899080834, - 0.016343594360),
    to_complex(0.011826304753, 0.004203947000),
    to_complex(- 0.008683879962, 0.009595157780),
    to_complex(0.006239196457, - 0.001581018480),
    to_complex(0.002213200462, 0.020197008950),
    to_complex(0.007159057738, - 0.005497735241),
    to_complex(- 0.014502753750, 0.024653659802),
    to_complex(- 0.010356255009, - 0.002071567732),
    to_complex(- 0.001934357810, 0.011846384408),
    to_complex(0.001354209876, - 0.004047522337),
    to_complex(- 0.006371757656, 0.029752846406),
    to_complex(0.004687542557, - 0.012038954146),
    to_complex(- 0.005339908826, 0.007900215132),
    to_complex(0.007712313608, 0.006390688550),
    to_complex(- 0.012688164516, 0.009224566157),
    to_complex(- 0.010908197879, 0.002402023381),
    to_complex(0.001505943505, 0.014791661906),
    to_complex(0.016891832491, 0.001316387415),
    to_complex(0.001616773027, 0.020638697927),
    to_complex(- 0.017960052425, 0.004544412412),
    to_complex(- 0.004747686337, - 0.008962016683),
    to_complex(- 0.002449902424, - 0.006527649144),
    to_complex(- 0.013365698875, 0.016015199813),
    to_complex(0.006137667728, - 0.010469210878),
    to_complex(0.000145709339, - 0.004114969359),
    to_complex(- 0.007935400320, 0.001080345126),
    to_complex(- 0.002228795123, 0.004116800778),
    to_complex(- 0.005112465838, 0.006909671552),
    to_complex(- 0.007182127344, 0.001861856952),
    to_complex(0.006395712345, - 0.002880648251),
    to_complex(- 0.010708571200, 0.012409929872),
    to_complex(- 0.003200802912, - 0.004772404873),
    to_complex(- 0.005184353441, 0.000590091092),
    to_complex(- 0.009347831423, 0.013251876980),
    to_complex(- 0.008252625250, - 0.003355245556),
    to_complex(- 0.004396822447, - 0.013712169332),
    to_complex(0.002949575420, - 0.001193337895),
    to_complex(0.007521208472, 0.005456543076),
    to_complex(- 0.007576470887, 0.010847848254),
    to_complex(- 0.001518611277, 0.002822546005),
    to_complex(- 0.002819677226, - 0.001262550660),
    to_complex(0.003755896210, - 0.006751239017),
    to_complex(- 0.013722387133, 0.010470010851),
    to_complex(0.001021040892, 0.005726781214),
    to_complex(- 0.000819185220, 0.005295596133),
    to_complex(0.001731111221, 0.002533886183),
    to_complex(0.001421904343, 0.005678943980),
    to_complex(- 0.011043514775, 0.001374994003),
    to_complex(0.005503252828, - 0.001308261496),
    to_complex(- 0.004646002490, - 0.004104029493),
    to_complex(- 0.001508599105, 0.007140897052),
    to_complex(- 0.004469113683, 0.014526115439),
    to_complex(- 0.003279041783, 0.009156784020),
    to_complex(0.007469025672, 0.005274507751),
    to_complex(0.003568155602, 0.020546963603),
    to_complex(0.000882469737, 0.000840861093),
    to_complex(0.001421122538, - 0.008525793023),
    to_complex(0.001839078176, - 0.005103582003),
    to_complex(- 0.016561775021, - 0.004071005999),
    to_complex(- 0.011318617577, - 0.003209579209),
    to_complex(0.007549911629, 0.004917941930),
    to_complex(0.001999451274, - 0.003607686227),
    to_complex(- 0.004711261955, 0.007442573155),
    to_complex(- 0.002778583699, 0.001455961555),
    to_complex(0.001275645168, - 0.004035469197),
    to_complex(0.001681769733, - 0.008403662214),
    to_complex(0.002016658814, 0.005979777607),
    to_complex(- 0.005511278134, 0.002545829154),
    to_complex(- 0.008734533656, - 0.007249735097),
    to_complex(0.007031159540, 0.003904248056),
    to_complex(0.007964029282, 0.013159687396),
    to_complex(- 0.006353880398, 0.006602783948),
    to_complex(0.006609563042, 0.000664163984),
    to_complex(0.001478509611, 0.007779941027),
    to_complex(- 0.002997080509, 0.007042970301),
    to_complex(0.000142769508, 0.006274122845),
    to_complex(- 0.003652354502, 0.002727145127),
    to_complex(0.006751795926, - 0.010786669180),
    to_complex(- 0.006862255137, 0.018632876683),
    to_complex(- 0.005082859459, - 0.001698961465),
    to_complex(0.001739538822, - 0.007365605422),
    to_complex(0.015463343741, 0.005046820013),
    to_complex(- 0.002515867773, 0.013902011991),
    to_complex(- 0.009255150170, 0.001632295297),
    to_complex(0.008712305411, - 0.003428344518),
    to_complex(0.001851072946, 0.005365830955),
    to_complex(0.002878237524, 0.001102978615),
    to_complex(- 0.005375291552, - 0.005131588375),
    to_complex(- 0.002485015338, 0.012435887936),
    to_complex(- 0.004589320347, - 0.001935004692),
    to_complex(0.002932091776, 0.019416569844),
    to_complex(0.000581733074, 0.001486896137),
    to_complex(- 0.007797724739, - 0.003902372431),
    to_complex(- 0.002038254345, - 0.001579579126),
    to_complex(0.000989769475, 0.010188405926),
    to_complex(- 0.008694273476, - 0.004213763260),
    to_complex(0.004499095849, 0.010435003465),
    to_complex(- 0.009252618978, - 0.005702114939),
    to_complex(0.003289095411, 0.002705889793),
    to_complex(- 0.005934878316, 0.002577413739),
    to_complex(- 0.002869506733, 0.003057351303),
    to_complex(0.009900424328, 0.009764051929),
    to_complex(- 0.007938403076, - 0.008381792380),
    to_complex(- 0.010354385360, - 0.001843919852),
    to_complex(0.010762644738, 0.002554923392),
    to_complex(- 0.003484904310, - 0.005965367764),
    to_complex(0.001824950458, 0.006049086071),
    to_complex(0.001840962134, 0.004416586202),
    to_complex(0.002195405953, 0.004431049707),
    to_complex(0.005673311561, 0.002563351659),
    to_complex(- 0.006127782304, - 0.000448713099),
    to_complex(0.004096522903, 0.003936962195),
    to_complex(0.005730664808, 0.001687285055),
    to_complex(0.005085719713, 0.012414620255),
    to_complex(- 0.016158464357, 0.014905276994),
    to_complex(- 0.006885285782, - 0.009781291330),
    to_complex(- 0.004021214343, 0.004504783063),
    to_complex(0.011885435414, - 0.000129555056),
    to_complex(0.005198134231, 0.009471465606),
    to_complex(- 0.005073927556, - 0.000219046566),
    to_complex(0.010837076214, - 0.001809889692),
    to_complex(0.003992937223, - 0.002469737677),
    to_complex(0.002701109128, 0.004137714771),
    to_complex(- 0.017953369337, - 0.012727488843),
    to_complex(- 0.004225761862, 0.005222136492),
    to_complex(- 0.002627140896, - 0.013331956475),
    to_complex(- 0.002625831943, 0.022111029500),
    to_complex(0.000044838170, - 0.004962879863),
    to_complex(0.000738763293, - 0.001552225686),
    to_complex(- 0.004438682729, - 0.002627432982),
    to_complex(0.010397618299, 0.012161743614),
    to_complex(0.002719219319, - 0.000591606559),
    to_complex(0.003568438527, - 0.009896095606),
    to_complex(0.011345019937, - 0.015990760524),
    to_complex(- 0.003545506030, 0.007870260535),
    to_complex(- 0.002492882066, - 0.001447333599),
    to_complex(0.010862701452, 0.010382072662),
    to_complex(0.011741598071, - 0.002594458503),
    to_complex(- 0.012270444126, 0.011423603073),
    to_complex(0.012490615451, 0.003949258618),
    to_complex(0.002396231104, - 0.010034152558),
    to_complex(- 0.001114604113, 0.005608767510),
    to_complex(- 0.003262005888, 0.008434488580),
    to_complex(- 0.005878375137, - 0.008948087939),
    to_complex(- 0.004157627245, - 0.000872820953),
    to_complex(0.009753039865, - 0.003092228911),
    to_complex(0.011615840986, 0.025174714714),
    to_complex(0.006598941643, - 0.002480132362),
    to_complex(0.004228235017, 0.004790393185),
    to_complex(0.008326205309, 0.008637567531),
    to_complex(- 0.007467354256, 0.019086720788),
    to_complex(0.009104710050, - 0.010863086253),
    to_complex(0.011778067992, - 0.004729880429),
    to_complex(- 0.007104621098, - 0.011631379351),
    to_complex(- 0.006551998392, 0.008666683476),
    to_complex(0.008784613472, 0.005711938613),
    to_complex(- 0.000785336220, 0.002110154289),
    to_complex(0.000203096027, - 0.007313178323),
    to_complex(- 0.017282280432, 0.022062593272),
    to_complex(- 0.002222496217, - 0.004635900072),
    to_complex(- 0.003431337295, 0.010107653074),
    to_complex(- 0.001329115876, 0.000373151148),
    to_complex(- 0.011879981700, 0.016080153061),
    to_complex(0.001500864803, 0.005267289684),
    to_complex(0.020157446151, 0.023364117670),
    to_complex(- 0.001525795751, 0.001273575272),
    to_complex(- 0.001571630235, 0.004275250318),
    to_complex(0.000727929682, 0.008712834963),
    to_complex(- 0.004945374762, - 0.002248738250),
    to_complex(0.006340463519, - 0.002572774405),
    to_complex(- 0.000826842467, 0.007104948578),
    to_complex(- 0.006224103960, - 0.001804787062),
    to_complex(- 0.000287389312, 0.002657789578),
    to_complex(0.007175238730, 0.006385992681),
    to_complex(- 0.007542451114, 0.001039415842),
    to_complex(- 0.001127494856, 0.005144987847),
    to_complex(0.000624300832, - 0.006483547471),
    to_complex(- 0.003472569057, - 0.005972554589),
    to_complex(0.007962343971, - 0.013639435910),
    to_complex(- 0.010956270358, 0.001148633459),
    to_complex(0.005382806365, 0.006370835744),
    to_complex(- 0.004034238703, 0.000765753464),
    to_complex(- 0.002310131373, 0.009387642265),
    to_complex(0.005642650052, - 0.000308464440),
    to_complex(0.002090843564, 0.005013500049),
    to_complex(- 0.010826053186, 0.005738012610),
    to_complex(- 0.006572080228, 0.010994649318),
    to_complex(- 0.008496746409, - 0.000172609428),
    to_complex(- 0.006467269112, - 0.010353221960),
    to_complex(0.005214287772, 0.004889941185),
    to_complex(0.000629861584, - 0.000968264895),
    to_complex(- 0.011501026029, - 0.004155521666),
    to_complex(0.023712545749, - 0.007398536503),
    to_complex(0.003017763038, 0.003979046296),
    to_complex(- 0.013928168182, - 0.000569710424),
    to_complex(- 0.003420223929, - 0.001711328964),
    to_complex(- 0.004212010578, 0.003251699253),
    to_complex(- 0.003595075811, 0.007366993016),
    to_complex(- 0.006771394797, 0.003770681423),
    to_complex(0.007014067146, 0.000786904134),
    to_complex(0.002591342417, - 0.004768799014),
    to_complex(0.002078241783, - 0.008635182332),
    to_complex(- 0.001468876883, 0.014109173240),
    to_complex(- 0.001746383007, 0.002730867499),
    to_complex(- 0.002883492877, 0.006332641883),
    to_complex(- 0.005159177593, - 0.004453182304),
    to_complex(- 0.013633207187, 0.015874529745),
    to_complex(- 0.000992794089, - 0.008438623826),
    to_complex(- 0.002997830044, 0.002338623808),
    to_complex(- 0.004171812183, 0.002866483201),
    to_complex(- 0.002514037873, - 0.003792315961),
    to_complex(0.000956954471, 0.005388150432),
    to_complex(0.000041406284, 0.011423883570),
    to_complex(0.007169625411, 0.008889455645),
    to_complex(0.003798594908, 0.008000010645),
    to_complex(0.003473625731, 0.001856179263),
    to_complex(0.001365547670, - 0.002387865219),
    to_complex(- 0.003299754474, - 0.006293720123),
    to_complex(0.014786547295, 0.003682926978),
    to_complex(0.009939587450, 0.002479223403),
    to_complex(- 0.008587121632, - 0.001538162773),
    to_complex(0.003424599693, 0.015322337437),
    to_complex(- 0.013048942928, 0.011252333939),
    to_complex(0.006304032945, 0.002776462119),
    to_complex(0.000447808559, - 0.001649438838),
    to_complex(- 0.004830419011, - 0.000443486948),
    to_complex(- 0.020821400202, 0.001569801823),
    to_complex(- 0.017900999362, 0.008920606913),
    to_complex(0.015021606905, - 0.007296941597),
    to_complex(- 0.010668982509, - 0.002657823868),
    to_complex(0.005077383983, 0.003454234550),
    to_complex(- 0.007062178909, 0.011209542682),
    to_complex(0.002463377250, 0.006268449261),
    to_complex(0.009868111476, - 0.001736246403),
    to_complex(0.004111487802, 0.007803709753),
    to_complex(0.006043124290, 0.002799370340),
    to_complex(0.002530661862, - 0.003555987536),
    to_complex(- 0.001160814714, - 0.005421004536),
    to_complex(0.014405385052, 0.014004101729),
    to_complex(0.006111371624, 0.003349306897),
    to_complex(- 0.009017433698, 0.003206270860),
    to_complex(- 0.006140332415, 0.008915184579),
    to_complex(0.005366345145, 0.000216744735),
    to_complex(0.000671350460, 0.004145641212),
    to_complex(0.001854184466, 0.008199893471),
    to_complex(0.003617458074, 0.010360630621),
    to_complex(- 0.004506673061, 0.009029063775),
    to_complex(0.000260789081, - 0.000674378381),
    to_complex(0.014249234986, 0.005241926315),
    to_complex(0.000763180903, - 0.005407310941),
    to_complex(- 0.008741808661, - 0.008415165621),
    to_complex(- 0.018651321440, 0.002993929848),
    to_complex(0.005263872044, - 0.002899261725),
    to_complex(0.002647982263, - 0.002002958352),
    to_complex(0.002263982608, 0.006535000959),
    to_complex(- 0.001638366459, 0.001232357073),
    to_complex(- 0.009447134175, 0.003437501276),
    to_complex(0.010144366677, - 0.007287034033),
    to_complex(0.014670335363, 0.005438051260),
    to_complex(0.000137647984, - 0.006327791548),
    to_complex(0.002939472008, 0.000596734542),
    to_complex(0.002825146025, - 0.007591393521),
    to_complex(0.003948577463, - 0.000211451773),
    to_complex(- 0.004197904415, - 0.003183282030),
    to_complex(- 0.007183872754, 0.000082863975),
    to_complex(0.005296243739, - 0.006766999599),
    to_complex(- 0.001012292395, 0.006442084876),
    to_complex(- 0.001146900078, - 0.003323422491),
    to_complex(- 0.009416702065, 0.005240545094),
    to_complex(0.008059742560, 0.004630189634),
    to_complex(0.001486375230, 0.016398188135),
    to_complex(- 0.005794841751, - 0.011325677844),
    to_complex(- 0.009892869553, - 0.010073558350),
    to_complex(0.005634409689, 0.013823070438),
    to_complex(0.000953703241, 0.003085534592),
    to_complex(0.002262335225, 0.000705029844),
    to_complex(0.001791310109, 0.004437492184),
    to_complex(0.012871591222, - 0.000659312177),
    to_complex(- 0.002029923384, - 0.003017497912),
    to_complex(- 0.004298401051, - 0.000424706270),
    to_complex(0.000646033465, - 0.003477719603),
    to_complex(0.012658939648, 0.013714541057),
    to_complex(- 0.001765702202, 0.019058106430),
    to_complex(- 0.001172935499, 0.002491530011),
    to_complex(0.001952756805, - 0.004283403980),
    to_complex(0.001419669917, 0.000633636394),
    to_complex(- 0.000138892162, 0.009121540757),
    to_complex(- 0.006560666484, - 0.007544244506),
    to_complex(- 0.005609624973, 0.006587068742),
    to_complex(- 0.001026074654, - 0.001314755089),
    to_complex(0.000253867920, - 0.002655545269),
    to_complex(0.001463597550, - 0.006948860147),
    to_complex(- 0.009594396977, 0.007902926644),
    to_complex(0.013252491094, - 0.000689492296),
    to_complex(- 0.001111122513, 0.017575006425),
    to_complex(- 0.002954422413, - 0.003128809642),
    to_complex(0.008925454501, 0.000598473650),
    to_complex(- 0.000340347413, - 0.014923822716),
    to_complex(0.004699079052, 0.009206892417),
    to_complex(- 0.006089145747, - 0.012015846776),
    to_complex(- 0.011160899591, - 0.007456957021),
    to_complex(0.002953728127, 0.002404749674),
    to_complex(- 0.001699102813, 0.018917312937),
    to_complex(0.004927403022, - 0.000975429025),
    to_complex(- 0.010146208167, - 0.000013574744),
    to_complex(0.008474271367, 0.008332751894),
    to_complex(- 0.002864579276, 0.008366693544),
    to_complex(0.003046504646, - 0.000556591035),
    to_complex(0.004422967048, - 0.001062361794),
    to_complex(0.003606286047, - 0.005179281344),
    to_complex(0.001007358402, 0.010397365476),
    to_complex(- 0.007388032759, - 0.001616266978),
    to_complex(0.005108932284, 0.000831763894),
    to_complex(0.003697926199, 0.010836187008),
    to_complex(0.010642527471, 0.000965268371),
    to_complex(- 0.004712612511, - 0.003752267435),
    to_complex(0.007308020891, 0.003094891374),
    to_complex(0.017401771771, 0.002778964030),
    to_complex(- 0.002052902121, 0.008866389361),
    to_complex(- 0.004956932764, 0.012785070654),
    to_complex(- 0.000507317719, - 0.006655345914),
    to_complex(0.001151848129, - 0.001858257858),
    to_complex(- 0.003951639565, 0.002838646681),
    to_complex(0.002112566618, - 0.005601978571),
    to_complex(- 0.000577098764, - 0.002708611957),
    to_complex(0.003903504733, 0.013176339542),
    to_complex(- 0.001678500870, 0.001638150036),
    to_complex(0.017239830925, 0.003232338789),
    to_complex(0.005690766946, - 0.008979755455),
    to_complex(0.006310646876, - 0.006344953466),
    to_complex(0.004800606391, 0.013307467863),
    to_complex(- 0.006385959668, - 0.003714597167),
    to_complex(0.004040720513, - 0.002265902593),
    to_complex(- 0.006525368486, - 0.004357622313),
    to_complex(0.014942231395, 0.014869855241),
    to_complex(0.004086713128, - 0.012317147944),
    to_complex(- 0.014812946893, 0.001572642474),
    to_complex(0.004663386906, - 0.004968130546),
    to_complex(- 0.001282031075, 0.010352962559),
    to_complex(0.001623745126, - 0.011282027323),
    to_complex(0.000443244777, 0.012712010701),
    to_complex(0.006716185455, - 0.003130232238),
    to_complex(0.001008242435, 0.021279863072),
    to_complex(- 0.007687874656, - 0.004512458725),
    to_complex(0.000079049215, - 0.006713223886),
    to_complex(0.008872514376, 0.001884624135),
    to_complex(0.000339562542, - 0.000266678035),
    to_complex(- 0.005384655360, 0.002389251193),
    to_complex(0.001634437639, 0.003125977466),
    to_complex(- 0.004556648323, 0.002740493338),
    to_complex(- 0.001923899720, 0.007487439727),
    to_complex(- 0.005010112707, - 0.000051141397),
    to_complex(- 0.003578224588, - 0.005348072134),
    to_complex(0.019530662484, - 0.004946559304),
    to_complex(0.016223138382, 0.018197790156),
    to_complex(- 0.009218171529, - 0.014649161729),
    to_complex(0.000099207041, - 0.006952200469),
    to_complex(- 0.003329422284, 0.001910523948),
    to_complex(0.015365169878, 0.009876560914),
    to_complex(0.012968418708, - 0.003277957280),
    to_complex(0.000833603752, 0.002010450027),
    to_complex(- 0.004530608724, - 0.002262294883),
    to_complex(- 0.000390043053, 0.013228326856),
    to_complex(0.006842352879, 0.003137187953),
    to_complex(0.004363166239, - 0.003603984173),
    to_complex(- 0.007872343721, - 0.016301604830),
    to_complex(0.003018002833, 0.009563727114),
    to_complex(0.002489384304, 0.014841780834),
    to_complex(0.006293984851, 0.003517762057),
    to_complex(- 0.005144024197, - 0.002416058831),
    to_complex(- 0.003486530856, 0.018204595651),
    to_complex(- 0.012743803704, 0.001256879384),
    to_complex(0.002411243638, 0.012193575594),
    to_complex(0.004324988622, 0.001666245027),
    to_complex(0.009299741787, 0.011365277028),
    to_complex(- 0.020388916154, 0.012004428525),
    to_complex(- 0.002044533159, 0.005485982461),
    to_complex(0.013803251013, 0.017111799353),
    to_complex(0.001607090631, - 0.002133716733),
    to_complex(- 0.003021931995, - 0.008588175451),
    to_complex(- 0.000978267303, 0.008568552828),
    to_complex(0.000057366187, - 0.003779354309),
    to_complex(0.002489772225, 0.006877297507),
    to_complex(- 0.000679961577, 0.007227438176),
    to_complex(- 0.007260640721, 0.002050949126),
    to_complex(0.006018101035, - 0.000858738177),
    to_complex(0.003198301487, 0.009548721049),
    to_complex(0.001520154010, - 0.006764964008),
    to_complex(- 0.007469920574, - 0.000338370547),
    to_complex(0.010466567400, 0.008508651966),
    to_complex(- 0.001753974126, 0.008849762787),
    to_complex(0.000873705308, 0.019351649883),
    to_complex(0.010789017579, 0.008564316245),
    to_complex(0.006825428417, 0.012005403333),
    to_complex(- 0.011054390206, 0.007969726754),
    to_complex(- 0.001450679493, - 0.008332268693),
    to_complex(0.001708859980, - 0.004740346960),
    to_complex(0.001675225163, 0.010368187030),
    to_complex(- 0.005803690725, - 0.000705069290),
    to_complex(0.001930837601, 0.006677276732),
    to_complex(- 0.002102030566, 0.004345130801),
    to_complex(0.000435741954, - 0.007366975033),
    to_complex(0.008480025275, 0.013212286678),
    to_complex(- 0.004938130746, - 0.008175388796),
    to_complex(- 0.003842401141, 0.001278555914),
    to_complex(- 0.003452630279, - 0.006626575853),
    to_complex(0.003282387887, 0.008249332875),
    to_complex(- 0.003428074901, - 0.000461361181),
    to_complex(- 0.015131483500, - 0.010442639166),
    to_complex(- 0.003283967996, 0.007157699615),
    to_complex(0.004587960473, 0.013993400342),
    to_complex(- 0.002279992569, 0.003404151696),
    to_complex(- 0.000200805596, - 0.002320562017),
    to_complex(0.017861611640, - 0.013768018033),
    to_complex(- 0.008722525237, 0.000084016848),
    to_complex(0.000201497340, 0.002521030555),
    to_complex(- 0.009372372145, 0.000908410222),
    to_complex(- 0.005666611623, - 0.000705579978),
    to_complex(0.001239671183, 0.007248626686),
    to_complex(- 0.009892708674, 0.008643179870),
    to_complex(- 0.000120919461, 0.006789072694),
    to_complex(0.004697587857, - 0.011945389284),
    to_complex(0.006505556300, 0.006188795460),
    to_complex(0.009960284170, - 0.013896963579),
    to_complex(- 0.003147655286, 0.014180181227),
    to_complex(0.006858708302, 0.010742862792),
    to_complex(- 0.006840005420, 0.015045567584),
    to_complex(0.004269161857, 0.002530711513),
    to_complex(- 0.000246938521, 0.005154133132),
    to_complex(0.000850609060, - 0.002944371875),
    to_complex(0.000088733425, 0.013228095614),
    to_complex(- 0.003197815945, - 0.002209631427),
    to_complex(0.005742344831, - 0.011102673959),
    to_complex(- 0.003874052863, 0.005977186697),
    to_complex(0.005720397052, 0.017513647532),
    to_complex(0.001771109998, 0.004481941229),
    to_complex(- 0.002119880650, - 0.018953650958),
    to_complex(- 0.008924289685, 0.006252252612),
    to_complex(0.003450762788, 0.022259441890),
    to_complex(0.011179094127, - 0.014164184191),
    to_complex(0.002853542026, 0.011080153494),
    to_complex(- 0.004646263096, 0.007236442384),
    to_complex(- 0.005320618418, - 0.000855262470),
    to_complex(- 0.004767559448, - 0.003916022059),
    to_complex(0.004956989118, - 0.016422467579),
    to_complex(0.008724933702, 0.017006034585),
    to_complex(0.000449217940, - 0.002189202544),
    to_complex(0.004680508566, 0.000636909508),
    to_complex(0.013700214502, - 0.002628064791),
    to_complex(0.002177816338, 0.001590981986),
    to_complex(0.005221923203, 0.006451741381),
    to_complex(0.012222303474, - 0.009469743279),
    to_complex(- 0.013603960091, - 0.000055475648),
    to_complex(- 0.000833012915, - 0.000466825068),
    to_complex(0.013213693140, 0.003241665686),
    to_complex(0.000124255604, 0.002560640581),
    to_complex(0.006466622811, - 0.005254577565),
    to_complex(- 0.006821955514, - 0.008986386595),
    to_complex(0.013282490387, 0.003475840460),
    to_complex(0.006121150226, - 0.004165026610),
    to_complex(0.007032559440, - 0.009193481592),
    to_complex(- 0.001967190890, 0.004562552945),
    to_complex(0.003642013856, 0.003534750896),
    to_complex(- 0.001717204177, 0.003971723141),
    to_complex(0.010033293396, - 0.002472330123),
    to_complex(- 0.006586896363, 0.002477366478),
    to_complex(0.001465866955, 0.010272008614),
    to_complex(- 0.013236239639, 0.000893282435),
    to_complex(0.002039358375, - 0.008683980005),
    to_complex(0.005605137647, - 0.002637886255),
    to_complex(- 0.002066079217, - 0.001411140586),
    to_complex(- 0.004124238614, 0.003945235500),
    to_complex(0.008851804006, - 0.002931935917),
    to_complex(- 0.000066499975, - 0.005626465430),
    to_complex(- 0.005885355165, 0.009921964804),
    to_complex(- 0.005469154344, 0.007039977720),
    to_complex(- 0.004508528973, - 0.008238334411),
    to_complex(0.005096108902, - 0.000665473471),
    to_complex(0.000706042931, 0.009488462574),
    to_complex(0.005470158741, - 0.000025803784),
    to_complex(- 0.001105222825, 0.013120990444),
    to_complex(0.000465613262, - 0.002421327949),
    to_complex(0.005023034435, 0.009967069240),
    to_complex(- 0.002606202118, - 0.008034043505),
    to_complex(- 0.002466016314, - 0.004934253919),
    to_complex(0.000178176371, 0.002576019716),
    to_complex(0.011378760043, 0.010320524869),
    to_complex(- 0.001381335317, 0.002615879335),
    to_complex(- 0.014559389890, 0.015356624117),
    to_complex(- 0.006412127542, - 0.004114654093),
    to_complex(0.002754558215, 0.001653945948),
    to_complex(0.008647436536, 0.007850822948),
    to_complex(- 0.015827698573, - 0.005804940471),
    to_complex(- 0.005508458251, 0.015127741368),
    to_complex(- 0.010856986485, 0.001675887856),
    to_complex(- 0.001587437265, - 0.001612625281),
    to_complex(- 0.002107765831, 0.007981841742),
    to_complex(0.007547135468, - 0.006096540831),
    to_complex(- 0.010827980538, 0.012221365523),
    to_complex(0.001469778292, 0.006157261268),
    to_complex(0.002202508999, - 0.007598209131),
    to_complex(0.011759714491, 0.005337622937),
    to_complex(0.004104819775, 0.007983175923),
    to_complex(0.000461642047, - 0.003367317420),
    to_complex(0.007015773714, - 0.004459445154),
    to_complex(0.001749362483, - 0.000432200057),
    to_complex(- 0.003914014682, 0.007259227469),
    to_complex(- 0.001918587913, - 0.005274112424),
    to_complex(- 0.001120728493, 0.002234042976),
    to_complex(- 0.012769982966, - 0.001444747150),
    to_complex(- 0.006682054678, - 0.000425589747),
    to_complex(0.000909777802, - 0.006619094642),
    to_complex(- 0.001662498134, - 0.003983609457),
    to_complex(- 0.007492878596, - 0.006272597219),
    to_complex(0.004394857868, 0.013065916486),
    to_complex(0.002025552571, - 0.007452941868),
    to_complex(0.006512232885, 0.000941895954),
    to_complex(0.002667399396, 0.003093087444),
    to_complex(0.007346110898, - 0.001396399638),
    to_complex(0.007163492704, 0.003198394763),
    to_complex(- 0.015968541034, - 0.003416021177),
    to_complex(0.009578092608, - 0.006838352615),
    to_complex(- 0.003903718042, - 0.004901646678),
    to_complex(0.000155631003, - 0.006116619298),
    to_complex(0.006762792747, 0.012130675012),
    to_complex(- 0.003710448749, - 0.011710224759),
    to_complex(0.005441012372, 0.000781304541),
    to_complex(0.002080750506, - 0.007561064964),
    to_complex(- 0.002386259770, 0.005383519196),
    to_complex(- 0.002430603363, - 0.007100142806),
    to_complex(- 0.005929209551, 0.002234547629),
    to_complex(0.006475732477, 0.005722016843),
    to_complex(0.000502591040, 0.006584659258),
    to_complex(0.002890049008, - 0.008342766051),
    to_complex(0.000220733494, 0.003988740217),
    to_complex(0.009782230018, 0.003293519130),
    to_complex(- 0.010906062974, - 0.000076083184),
    to_complex(- 0.008382972583, 0.012592457416),
    to_complex(0.011087389994, 0.014474145195),
    to_complex(- 0.011551989708, 0.010052048908),
    to_complex(- 0.012196096986, - 0.014524061575),
    to_complex(0.007008301834, - 0.003115432183),
    to_complex(0.006634266480, 0.003596270945),
    to_complex(- 0.001957556762, - 0.007051916590),
    to_complex(- 0.004999748347, - 0.005588630498),
    to_complex(- 0.005323103459, 0.004494628174),
    to_complex(- 0.002587748265, - 0.004615656820),
    to_complex(- 0.001676427928, 0.008915158597),
    to_complex(0.003807067789, 0.011761450808),
    to_complex(- 0.002667215530, - 0.000548924231),
    to_complex(- 0.008767358851, 0.017950064326),
    to_complex(- 0.001118853297, 0.012008673742),
    to_complex(- 0.005196225322, 0.000557188776),
    to_complex(0.003510268871, - 0.003478292529),
    to_complex(- 0.012970428886, 0.011235321397),
    to_complex(- 0.007067859375, - 0.004045956660),
    to_complex(0.003461212160, - 0.001246804827),
    to_complex(- 0.005536831694, 0.007833919525),
    to_complex(0.012736530430, - 0.001962334836),
    to_complex(0.003975699171, - 0.004272708859),
    to_complex(- 0.005848734256, 0.006207006434),
    to_complex(0.002080247101, - 0.013658308353),
    to_complex(0.002406202103, 0.011738015479),
    to_complex(- 0.010708342080, - 0.000008206011),
    to_complex(0.001187837282, - 0.001045766145),
    to_complex(0.004179888450, - 0.001756921054),
    to_complex(0.011535422702, 0.002388968076),
    to_complex(0.005652899631, 0.000278363461),
    to_complex(- 0.012115187791, - 0.003271252641),
    to_complex(0.005115593757, - 0.006252728412),
    to_complex(0.010789634369, 0.012242969585),
    to_complex(- 0.004563095405, 0.000655028829),
    to_complex(- 0.005600446834, 0.003231386415),
    to_complex(0.004117802814, 0.003313404131),
    to_complex(0.000953411695, 0.003855009694),
    to_complex(- 0.004341302925, - 0.001852491856),
    to_complex(- 0.002347895939, 0.003047483775),
    to_complex(- 0.001916967696, - 0.002832386409),
    to_complex(- 0.012117561533, 0.008719207898),
    to_complex(- 0.008921089849, - 0.007010377973),
    to_complex(0.003115751131, 0.000205365305),
    to_complex(0.001398583952, 0.000148696537),
    to_complex(0.008279396360, 0.014780118964),
    to_complex(- 0.017039691844, 0.013059100261),
    to_complex(0.012072080854, - 0.001601821533),
    to_complex(- 0.006404022460, - 0.005452987330),
    to_complex(0.006422418722, - 0.002391719792),
    to_complex(- 0.003456747127, - 0.003362447567),
    to_complex(- 0.001794766993, 0.000018224726),
    to_complex(0.010559280680, - 0.009521599749),
    to_complex(0.003921250163, 0.001600565046),
    to_complex(- 0.002187420386, 0.004608946729),
    to_complex(- 0.016157606788, 0.010075512571),
    to_complex(- 0.000656597615, 0.006228935566),
    to_complex(- 0.006197778537, 0.000459468464),
    to_complex(- 0.003587346696, - 0.013418214669),
    to_complex(- 0.007394654692, - 0.002816316324),
    to_complex(0.003876484088, 0.001749067158),
    to_complex(0.001145698657, 0.005277399041),
    to_complex(- 0.010552541588, - 0.003555122636),
    to_complex(- 0.003137008237, - 0.003981836819),
    to_complex(0.003561976601, 0.002405819321),
    to_complex(0.000778454003, 0.014690259738),
    to_complex(- 0.008063384387, 0.005162070547),
    to_complex(0.003767411232, - 0.015489440915),
    to_complex(0.004018928377, - 0.006681673352),
    to_complex(- 0.002577757802, - 0.002750197316),
    to_complex(- 0.002397770500, - 0.005681887565),
    to_complex(- 0.003599477739, 0.009799095284),
    to_complex(- 0.005378314314, 0.001826537101),
    to_complex(- 0.002940447740, 0.005015942496),
    to_complex(- 0.015501453906, - 0.000101042546),
    to_complex(0.002735686555, - 0.013434710763),
    to_complex(0.021456671780, - 0.002829146511),
    to_complex(0.005211474164, 0.000508601200),
    to_complex(0.003851530059, - 0.000406759742),
    to_complex(0.010261135959, - 0.005629968429),
    to_complex(- 0.007075738216, 0.003928592221),
    to_complex(- 0.001277687876, 0.002485321147),
    to_complex(- 0.015077364264, 0.002534073320),
    to_complex(0.005344372953, 0.004090059678),
    to_complex(- 0.003055755671, - 0.000527305832),
    to_complex(0.002650471771, 0.004986211281),
    to_complex(- 0.016560940939, 0.007214164857),
    to_complex(0.010227441786, 0.006571082140),
    to_complex(0.006711733748, - 0.009705600567),
    to_complex(- 0.000375189166, - 0.004247665589),
    to_complex(0.019094583565, 0.010378647136),
    to_complex(- 0.009676825572, - 0.001961379071),
    to_complex(- 0.008096070980, 0.000414332584),
    to_complex(0.008455783529, 0.006347584670),
    to_complex(0.005139636706, - 0.000943300885),
    to_complex(- 0.003896689923, 0.000927608260),
    to_complex(- 0.001152334327, - 0.003548743218),
    to_complex(- 0.000016047239, 0.012319291761),
    to_complex(- 0.005277192693, 0.004811277687),
    to_complex(- 0.002486515097, - 0.005361127112),
    to_complex(- 0.000418769647, 0.003907724292),
    to_complex(0.008091521743, - 0.004604493906),
    to_complex(0.005540387038, - 0.007458163785),
    to_complex(0.001712769557, - 0.008497957174),
    to_complex(0.001872147894, - 0.002246766964),
    to_complex(- 0.001755992326, 0.008176099021),
    to_complex(- 0.011121104295, 0.007336353191),
    to_complex(- 0.001273418616, - 0.004059592248),
    to_complex(- 0.005329949920, - 0.006490142749),
    to_complex(- 0.006894971508, 0.005854822832),
    to_complex(0.007933309041, 0.005325978097),
    to_complex(0.002925343704, - 0.008050130491),
    to_complex(0.014172516173, - 0.003726737250),
    to_complex(0.011593580957, 0.005171840256),
    to_complex(- 0.006508759415, - 0.002338173585),
    to_complex(- 0.009523014564, - 0.001671453308),
    to_complex(- 0.006971394285, - 0.004504341962),
    to_complex(- 0.002119887313, 0.016145021991),
    to_complex(- 0.012234606730, - 0.012047211615),
    to_complex(0.000424714896, 0.000724238015),
    to_complex(- 0.006706380467, 0.011768167987),
    to_complex(- 0.006411065133, 0.002071714556),
    to_complex(0.001050945068, 0.002270041404),
    to_complex(0.003031057781, - 0.014290879210),
    to_complex(0.002154564243, - 0.012301460783),
    to_complex(0.010216293917, - 0.005900103604),
    to_complex(0.001402557776, 0.011903487963),
    to_complex(0.001337965289, 0.005463279156),
    to_complex(- 0.007056927594, - 0.004524711963),
    to_complex(- 0.005651066464, 0.006339741618),
    to_complex(- 0.004214106770, 0.014286722080),
    to_complex(0.003994606891, - 0.006118939761),
    to_complex(0.002029178727, 0.002544410841),
    to_complex(0.006430714684, 0.010225817071),
    to_complex(- 0.001197056831, - 0.007830276183),
    to_complex(0.008385825456, - 0.008665992820),
    to_complex(- 0.008822210436, 0.001601587380),
    to_complex(0.024916964306, 0.008743438684),
    to_complex(- 0.000477784946, - 0.009268475889),
    to_complex(- 0.006366246386, 0.007595566167),
    to_complex(- 0.002669532723, - 0.003847619810),
    to_complex(- 0.017568314020, - 0.008572266724),
    to_complex(0.005301115909, 0.002446060214),
    to_complex(0.003230346219, 0.009147369825),
    to_complex(0.003442074267, - 0.002725001603),
    to_complex(0.016610247346, 0.014339231316),
    to_complex(0.004345215121, 0.006162962228),
    to_complex(0.013651040462, - 0.009596531310),
    to_complex(0.004743789683, - 0.006843539357),
    to_complex(0.010288974833, 0.004054665493),
    to_complex(0.009027682861, 0.009309956925),
    to_complex(0.006686318651, 0.003608688674),
    to_complex(- 0.000947713022, - 0.010745916674),
    to_complex(0.004532254748, 0.014107317912),
    to_complex(- 0.005431628386, 0.002229373129),
    to_complex(- 0.005157661269, 0.006128037090),
    to_complex(- 0.007905478499, - 0.005011313677),
    to_complex(0.001353701152, - 0.002832423134),
    to_complex(- 0.000266831837, - 0.006015664502),
    to_complex(- 0.011711320167, 0.007686574812),
    to_complex(0.002264551747, - 0.015223109938),
    to_complex(0.004695782655, 0.004469382085),
    to_complex(0.000134984764, - 0.003227081746),
    to_complex(0.003878431606, - 0.003176352122),
    to_complex(- 0.009634814838, - 0.004940820847),
    to_complex(- 0.007144021596, 0.002309011084),
    to_complex(0.003088873267, 0.002601226926),
    to_complex(- 0.011090295562, - 0.005070565446),
    to_complex(0.000674305381, - 0.007535155849),
    to_complex(0.005895826407, - 0.006274184101),
    to_complex(- 0.005298799924, - 0.006710721902),
    to_complex(- 0.003918102935, 0.009487611015),
    to_complex(0.012542402943, - 0.004078480911),
    to_complex(- 0.004876933769, - 0.006985276964),
    to_complex(0.006741048144, - 0.005367007018),
    to_complex(0.007381357802, 0.002162355032),
    to_complex(- 0.007382440735, - 0.001696051138),
    to_complex(- 0.006091723632, 0.004680240326),
    to_complex(0.003321302859, - 0.001589254795),
    to_complex(- 0.006649877650, 0.009404677755),
    to_complex(0.003955385893, - 0.005948365224),
    to_complex(0.002301943526, - 0.001474760894),
    to_complex(0.007025760876, - 0.012208331140),
    to_complex(0.007674921174, - 0.001098288185),
    to_complex(0.001891443603, - 0.003288426668),
    to_complex(0.012710020917, 0.007979525527),
    to_complex(- 0.005447658328, - 0.003020109320),
    to_complex(0.007142584503, - 0.008220906827),
    to_complex(- 0.011423311709, - 0.014871541657),
    to_complex(0.006244061898, 0.024299552641),
    to_complex(- 0.002263397411, 0.003620188467),
    to_complex(0.003098067351, 0.014482310721),
    to_complex(0.002418678629, 0.001980191500),
    to_complex(0.001571543527, - 0.006246237723),
    to_complex(- 0.010249471639, 0.007965997889),
    to_complex(- 0.004205643479, - 0.002974381921),
    to_complex(- 0.003670303120, 0.007667652372),
    to_complex(- 0.000602539977, 0.011368021712),
    to_complex(- 0.002538059641, 0.005651454721),
    to_complex(- 0.001676482958, 0.002489715477),
    to_complex(- 0.003793182801, - 0.002379402764),
    to_complex(0.013452932120, 0.017044845043),
    to_complex(- 0.005116194471, 0.000000221523),
    to_complex(- 0.009671910393, - 0.008642380842),
    to_complex(- 0.000379821466, - 0.009879679907),
    to_complex(0.016965688775, 0.005062654366),
    to_complex(- 0.015034826008, - 0.004853562666),
    to_complex(- 0.005466371237, - 0.011393825394),
    to_complex(- 0.004493624666, - 0.003335688745),
    to_complex(- 0.010127089096, 0.008543359433),
    to_complex(- 0.005104870315, 0.007769475413),
    to_complex(0.002322591107, - 0.000562225652),
    to_complex(0.012435608240, - 0.006115496572),
    to_complex(0.001273331885, 0.000476050409),
    to_complex(- 0.002394867934, - 0.009526676559),
    to_complex(0.007430579699, 0.001554486675),
    to_complex(0.002221796801, - 0.006414382302),
    to_complex(0.006046492559, - 0.000538987897),
    to_complex(- 0.003718135587, - 0.002398632249),
    to_complex(0.014394780735, - 0.001935720377),
    to_complex(0.013612104737, 0.001660393077),
    to_complex(- 0.004507028967, 0.003573343196),
    to_complex(- 0.002582137993, 0.009590189383),
    to_complex(- 0.001832767211, - 0.002752599972),
    to_complex(0.007795673700, 0.002897386333),
    to_complex(0.000147487006, - 0.004037921035),
    to_complex(0.003717154343, - 0.007529367349),
    to_complex(- 0.009240601256, - 0.013527810698),
    to_complex(0.001478629272, - 0.004764235563),
    to_complex(0.006769010425, 0.003492193115),
    to_complex(- 0.010103410990, - 0.000835794708),
    to_complex(- 0.003230037208, 0.002496947356),
    to_complex(0.007677185860, 0.000963147169),
    to_complex(0.018892900491, - 0.003684147738),
    to_complex(0.002064843150, 0.012374066803),
    to_complex(0.001348030895, 0.007593279978),
    to_complex(0.010893912180, 0.004008408661),
    to_complex(0.006364180652, 0.001177010645),
    to_complex(- 0.006887373824, 0.011212688627),
    to_complex(- 0.001081927910, 0.004793731592),
    to_complex(- 0.006948419433, 0.007217024538),
    to_complex(0.007168441861, - 0.001469256922),
    to_complex(0.003243808721, 0.009565586302),
    to_complex(- 0.004338062276, - 0.001365656915),
    to_complex(- 0.004364157024, - 0.006062646685),
    to_complex(0.011692159102, - 0.003346093203),
    to_complex(- 0.016447485931, - 0.004105659601),
    to_complex(0.006287000983, - 0.011371850073),
    to_complex(- 0.004163926829, - 0.005306481906),
    to_complex(0.016669310872, - 0.003012302189),
    to_complex(0.003588021752, 0.007354477840),
    to_complex(- 0.007222869069, 0.010774784575),
    to_complex(- 0.005543351991, - 0.004757027656),
    to_complex(0.009862947773, 0.002776067212),
    to_complex(- 0.010164991634, - 0.005582814256),
    to_complex(0.002103846951, 0.007334301368),
    to_complex(0.001057520621, - 0.010680271474),
    to_complex(- 0.004653634950, 0.013430767295),
    to_complex(0.003767174767, 0.005592763258),
    to_complex(- 0.001451707015, - 0.013497180085),
    to_complex(0.000717987625, - 0.004910448806),
    to_complex(0.003763394642, 0.000819082577),
    to_complex(0.004347057029, 0.004742066845),
    to_complex(- 0.001541393868, 0.008762894864),
    to_complex(0.007390970101, - 0.001515173703),
    to_complex(- 0.004329717195, - 0.000372385072),
    to_complex(- 0.000946505829, - 0.017304972955),
    to_complex(- 0.007654746591, - 0.004328226707),
    to_complex(- 0.009211330410, 0.006850904535),
    to_complex(0.008784111353, - 0.001564312819),
    to_complex(0.012897475815, 0.005197947993),
    to_complex(0.002579985731, 0.002686162106),
    to_complex(- 0.002632332359, - 0.011913580797),
    to_complex(0.005602258631, 0.001938985113),
    to_complex(- 0.001736707657, 0.007007457396),
    to_complex(0.009136129006, 0.003406742504),
    to_complex(0.004702948428, 0.003463362831),
    to_complex(0.005489429694, 0.003962776303),
    to_complex(0.007029798533, - 0.005544888559),
    to_complex(0.011937373116, 0.003340716850),
    to_complex(0.003047225664, 0.000253572182),
    to_complex(- 0.000414089696, 0.001584536412),
    to_complex(0.009546125005, - 0.009831788422),
    to_complex(0.001240868028, 0.000168173998),
    to_complex(0.005892954096, - 0.007109611100),
    to_complex(0.011486058764, 0.015003689886),
    to_complex(- 0.004484739514, 0.004298321448),
    to_complex(- 0.009314836285, 0.012784483857),
    to_complex(- 0.000959525813, - 0.000316561949),
    to_complex(0.015696634535, 0.001520065289),
    to_complex(- 0.003104334559, - 0.003076488604),
    to_complex(- 0.001281054545, - 0.004072956831),
    to_complex(- 0.005507051389, - 0.003875797993),
    to_complex(0.010963952082, 0.013397364656),
    to_complex(- 0.002169200746, - 0.007079318263),
    to_complex(- 0.006823774393, 0.005096744321),
    to_complex(0.000223343997, - 0.001851860618),
    to_complex(- 0.008961742986, 0.014040208169),
    to_complex(- 0.004393652138, - 0.008562927397),
    to_complex(0.000542976270, 0.002192346455),
    to_complex(0.000541684818, - 0.008339670680),
    to_complex(0.011170689317, - 0.000290505896),
    to_complex(- 0.009708677241, 0.000861896191),
    to_complex(0.000220781344, - 0.003509970658),
    to_complex(0.004585321638, 0.001486282096),
    to_complex(0.006821586882, 0.003549037470),
    to_complex(0.002341438474, 0.003387366104),
    to_complex(0.002211649894, - 0.010286777338),
    to_complex(0.001957044388, - 0.003593962952),
    to_complex(- 0.005558543889, - 0.000286335853),
    to_complex(- 0.001925280725, 0.000860102877),
    to_complex(- 0.000080233717, - 0.000464169427),
    to_complex(0.007911882328, 0.004627065477),
    to_complex(0.004766653699, 0.004242702967),
    to_complex(- 0.005238184720, 0.009684543493),
    to_complex(- 0.000484075644, 0.008178660625),
    to_complex(- 0.004278584591, - 0.011119826205),
    to_complex(0.005717766248, - 0.004849957276),
    to_complex(- 0.003391129851, - 0.004659987403),
    to_complex(0.000574164473, 0.001235154070),
    to_complex(0.005036339208, - 0.009663904320),
    to_complex(- 0.005160707256, 0.004999166801),
    to_complex(- 0.002525248735, 0.003877418001),
    to_complex(- 0.006778958389, - 0.001044704443),
    to_complex(0.001409691062, - 0.004097499006),
    to_complex(0.005994562037, 0.014996954287),
    to_complex(- 0.003013053483, - 0.000835961049),
    to_complex(0.010184158355, 0.004995399504),
    to_complex(0.006250061819, - 0.004971474877),
    to_complex(0.013559513041, 0.011833906642),
    to_complex(0.006093945609, - 0.012371923242),
    to_complex(0.013059961579, - 0.003612033095),
    to_complex(0.004736067307, - 0.001110610862),
    to_complex(0.008942625668, - 0.010825085978),
    to_complex(- 0.003393153059, 0.023000350793),
    to_complex(- 0.009804959856, - 0.001556828968),
    to_complex(- 0.003070393596, 0.014532749155),
    to_complex(0.007305540658, 0.007856596758),
    to_complex(0.005240067477, 0.000405235095),
    to_complex(- 0.005493190683, - 0.010465194523),
    to_complex(- 0.013287715863, - 0.004902638260),
    to_complex(0.008060241069, 0.004912609141),
    to_complex(0.005092844760, - 0.013191750585),
    to_complex(- 0.003948522298, - 0.004023680099),
    to_complex(0.006941988030, 0.002976667035),
    to_complex(0.002952976539, 0.008737012571),
    to_complex(0.002590054566, 0.000285488930),
    to_complex(0.001608122909, - 0.008601463495),
    to_complex(- 0.002726160556, - 0.010601894907),
    to_complex(- 0.001922657215, 0.003523976465),
    to_complex(- 0.005536191397, 0.002250269657),
    to_complex(0.010478605185, 0.012635669484),
    to_complex(- 0.008413830882, 0.002041429768),
    to_complex(0.008690654646, 0.003407939944),
    to_complex(- 0.003197628241, 0.001923070985),
    to_complex(0.000453633471, - 0.001789498328),
    to_complex(- 0.004141956592, - 0.005617784677),
    to_complex(0.011265723318, 0.009763804240),
    to_complex(- 0.002881595995, - 0.000099920667),
    to_complex(- 0.003442480161, 0.001810724589),
    to_complex(- 0.004737496132, 0.001179891069),
    to_complex(0.004132940808, - 0.003107783034),
    to_complex(0.002845542467, - 0.006019921427),
    to_complex(- 0.000292781046, - 0.003865594247),
    to_complex(0.012122537496, - 0.016561684787),
    to_complex(0.004472237023, 0.007249205283),
    to_complex(- 0.007305825571, 0.006796998829),
    to_complex(- 0.007218722261, 0.009430896574),
    to_complex(0.002355572249, - 0.012466101142),
    to_complex(0.013671869423, 0.011304349760),
    to_complex(0.001574723649, - 0.009287098777),
    to_complex(0.001811836940, - 0.004593287506),
    to_complex(0.002364417125, - 0.002757501037),
    to_complex(0.006130564874, - 0.009000546582),
    to_complex(- 0.006683711729, 0.004923837205),
    to_complex(- 0.003597145781, 0.000025506956),
    to_complex(0.002965705522, - 0.001831904190),
    to_complex(0.018666603593, - 0.007554734376),
    to_complex(0.006133733714, 0.004681085355),
    to_complex(0.007438472746, - 0.002957464588),
    to_complex(0.005989065984, 0.009118864717),
    to_complex(- 0.005116692890, 0.012764955436),
    to_complex(0.007503114066, 0.000306046589),
    to_complex(- 0.019296772633, 0.001315097402),
    to_complex(- 0.001720781558, 0.007179014213),
    to_complex(0.009126042304, 0.012303608676),
    to_complex(0.000623239621, 0.001945209777),
    to_complex(0.003465355477, 0.016490755321),
    to_complex(- 0.006544051565, 0.004675990384),
    to_complex(- 0.003063891182, 0.012128141087),
    to_complex(- 0.000744674528, - 0.002039338357),
    to_complex(- 0.002763327981, - 0.010130709310),
    to_complex(- 0.007510513135, 0.006408448881),
    to_complex(- 0.000914365601, 0.007221045778),
    to_complex(0.000346841605, 0.006293801714),
    to_complex(- 0.014402858579, - 0.005815202274),
    to_complex(- 0.010068321071, - 0.005558036873),
    to_complex(0.012352487198, 0.010655075003),
    to_complex(- 0.000505764755, - 0.001663242257),
    to_complex(0.017425789232, 0.010921867371),
    to_complex(0.003869786000, - 0.006788704991),
    to_complex(0.009787974733, 0.016606113704),
    to_complex(- 0.006158123722, - 0.011019208046),
    to_complex(0.010807816375, - 0.017236971582),
    to_complex(- 0.000293834361, 0.000234638465),
    to_complex(- 0.007031438626, 0.015704963080),
    to_complex(- 0.012106087011, 0.008518137515),
    to_complex(- 0.003810852249, 0.007889783924),
    to_complex(0.002720592776, - 0.002823777113),
    to_complex(- 0.011142073521, 0.004165593113),
    to_complex(- 0.006160116430, 0.003318851042),
    to_complex(- 0.002964240733, - 0.008734234923),
    to_complex(0.005165727991, 0.010199484853),
    to_complex(0.003377621126, 0.000076152678),
    to_complex(- 0.011478513528, 0.004559665783),
    to_complex(0.000692041673, - 0.002460388499),
    to_complex(0.016009505053, 0.011856737970),
    to_complex(0.002741455166, 0.013546564238),
    to_complex(- 0.000145393403, 0.006358953964),
    to_complex(0.006372721000, - 0.002781201919),
    to_complex(- 0.007035676425, - 0.010311666032),
    to_complex(- 0.012264184838, 0.004839147248),
    to_complex(0.005173380118, 0.009294563407),
    to_complex(- 0.003915993098, - 0.000955156211),
    to_complex(0.013920852725, - 0.011587027306),
    to_complex(- 0.001937606599, 0.016965323231),
    to_complex(- 0.001605922455, - 0.007571459798),
    to_complex(- 0.010828877664, 0.011269765598),
    to_complex(- 0.003885366451, 0.004116082394),
    to_complex(0.005916493793, 0.004479871843),
    to_complex(- 0.004035627185, 0.002101263152),
    to_complex(0.008591246064, 0.002882852456),
    to_complex(0.001027374623, - 0.004246411506),
    to_complex(0.000802084131, 0.006348968142),
    to_complex(0.006558597400, 0.005139819716),
    to_complex(- 0.014200839292, 0.006476005023),
    to_complex(0.000962310946, - 0.008880600318),
    to_complex(0.009139793213, 0.004284081291),
    to_complex(0.003894782391, 0.000374033690),
    to_complex(0.004939930117, 0.013584283688),
    to_complex(- 0.000262202403, - 0.013782567269),
    to_complex(0.011945886292, 0.007219278103),
    to_complex(- 0.000734460999, - 0.002751208887),
    to_complex(- 0.013828189167, - 0.007445120892),
    to_complex(- 0.000148298114, 0.007959663464),
    to_complex(- 0.000324352731, 0.009265409036),
    to_complex(- 0.007312054391, 0.007553099081),
    to_complex(- 0.002656129567, 0.015576792357),
    to_complex(- 0.004845656173, 0.003484662570),
    to_complex(0.003870313535, - 0.006013135369),
    to_complex(0.008851022780, 0.001167149641),
    to_complex(0.008616080759, - 0.007235407047),
    to_complex(0.011789008711, 0.001014201209),
    to_complex(0.000783687549, 0.001850006184),
    to_complex(0.001333848975, 0.005249998624),
    to_complex(0.013942420094, 0.005561787794),
    to_complex(0.004672805393, 0.010128204952),
    to_complex(- 0.001803983888, - 0.001426985308),
    to_complex(0.004698594467, 0.006081859573),
    to_complex(0.006787198374, - 0.007924585799),
    to_complex(- 0.001989490397, 0.006098402651),
    to_complex(0.000273373597, 0.009305533305),
    to_complex(0.001992841155, - 0.004002910030),
    to_complex(0.005329086806, 0.000019873309),
    to_complex(0.003853805356, 0.012042373437),
    to_complex(- 0.005833748070, - 0.007769328552),
    to_complex(- 0.002549558143, 0.003585627538),
    to_complex(- 0.009896056006, - 0.007028220252),
    to_complex(- 0.008353182642, - 0.007482230282),
    to_complex(0.010777764319, 0.008466012791),
    to_complex(- 0.001734838545, 0.005133179081),
    to_complex(0.000756541970, 0.007321002697),
    to_complex(- 0.003725774951, 0.008513438608),
    to_complex(0.012877394210, - 0.006712579607),
    to_complex(- 0.006900581856, - 0.004230713738),
    to_complex(- 0.013007955205, - 0.006824604326),
    to_complex(0.003457509561, - 0.000209915698),
    to_complex(0.008863992486, 0.012948911605),
    to_complex(- 0.000841221382, 0.002226834368),
    to_complex(0.015849675437, - 0.002529731251),
    to_complex(0.000735696577, - 0.000390573067),
    to_complex(0.002568767251, - 0.007243230705),
    to_complex(0.000348114209, - 0.004248983846),
    to_complex(- 0.003192412979, 0.000440351167),
    to_complex(0.008723647728, - 0.009152441962),
    to_complex(- 0.004999408161, - 0.006450102781),
    to_complex(- 0.008440438083, 0.017015410598),
    to_complex(- 0.000550126309, 0.004513744061),
    to_complex(- 0.003790654913, - 0.008037228738),
    to_complex(0.004050525470, - 0.004348138360),
    to_complex(- 0.000615741408, - 0.001377948726),
    to_complex(0.009532274029, - 0.005970805935),
    to_complex(0.005643500297, - 0.009717982124),
    to_complex(- 0.003097438181, 0.013897107477),
    to_complex(- 0.007714588156, 0.005981436717),
    to_complex(- 0.002494353747, 0.001046023307),
    to_complex(0.015182422787, 0.000231904293),
    to_complex(0.000329116416, - 0.004717149175),
    to_complex(- 0.004123555201, - 0.003290904095),
    to_complex(- 0.003446366018, 0.001076686919),
    to_complex(- 0.000994213179, - 0.007735154897),
    to_complex(- 0.011347890849, 0.009695733113),
    to_complex(0.005004072798, - 0.008667132113),
    to_complex(- 0.007619486954, 0.004691239244),
    to_complex(0.008065900158, - 0.005552599779),
    to_complex(0.013961402360, 0.011050996969),
    to_complex(- 0.013563743955, 0.004817844794),
    to_complex(0.008971942924, - 0.005398086833),
    to_complex(- 0.007534270513, - 0.002200214444),
    to_complex(- 0.003681506640, 0.002879599637),
    to_complex(- 0.003213208941, 0.007305268219),
    to_complex(- 0.006760052257, - 0.004999030761),
    to_complex(- 0.012154563710, 0.002913212266),
    to_complex(0.009881477834, - 0.000368465680),
    to_complex(0.004684934252, 0.006664614833),
    to_complex(0.002893632994, 0.006767042965),
    to_complex(- 0.002798909527, 0.012095614940),
    to_complex(0.011631445410, - 0.004190529107),
    to_complex(0.002165402698, - 0.002832541538),
    to_complex(- 0.005120260214, 0.013866063955),
    to_complex(0.004837155984, - 0.006715484138),
    to_complex(- 0.000736721612, 0.002013699219),
    to_complex(- 0.009880666088, - 0.000064821299),
    to_complex(0.000324984640, 0.007811512148),
    to_complex(0.002520881692, 0.001958313053),
    to_complex(- 0.003262156364, - 0.015716056320),
    to_complex(0.011326172090, 0.010598376860),
    to_complex(- 0.002636306586, - 0.010185112662),
    to_complex(0.006398058982, - 0.000510674906),
    to_complex(0.005219376076, 0.004311228033),
    to_complex(- 0.014955361431, 0.004969414929),
    to_complex(- 0.012440093812, 0.010295427208),
    to_complex(0.008389657991, - 0.013701701811),
    to_complex(- 0.001258379029, 0.006165027787),
    to_complex(0.016212787570, 0.006333573359),
    to_complex(- 0.000015634746, 0.012199604466),
    to_complex(0.007314105870, - 0.005229448038),
    to_complex(0.003366028093, - 0.004189604398),
    to_complex(- 0.005856106310, - 0.003056707918),
    to_complex(0.007891896591, - 0.002437548342),
    to_complex(- 0.005512112522, 0.006110830150),
    to_complex(- 0.007374117723, 0.001072558415),
    to_complex(- 0.011746350847, - 0.002031422807),
    to_complex(0.006575788921, - 0.000342840686),
    to_complex(- 0.002178266080, - 0.006677385137),
    to_complex(0.009469915270, 0.001349498098),
    to_complex(0.002853841091, 0.008028941485),
    to_complex(- 0.006354415263, - 0.005203062301),
    to_complex(0.001206899198, - 0.008286702884),
    to_complex(0.011418369209, 0.006693674954),
    to_complex(- 0.001345680959, - 0.000933096368),
    to_complex(0.001534733907, 0.002303893770),
    to_complex(- 0.000359815685, 0.008705270917),
    to_complex(0.012511513483, 0.003776964447),
    to_complex(- 0.007922452013, - 0.009468756562),
    to_complex(0.006939991876, - 0.014089952704),
    to_complex(- 0.006656728073, - 0.008981449875),
    to_complex(0.000980064280, 0.003309399028),
    to_complex(- 0.000011982538, - 0.004439326687),
    to_complex(- 0.005771121020, - 0.007149692616),
    to_complex(0.003589740564, - 0.001537308304),
    to_complex(0.011781991613, 0.002770949458),
    to_complex(0.010654841363, 0.014707059965),
    to_complex(0.007444753095, 0.001101023525),
    to_complex(0.005753404117, - 0.003663105557),
    to_complex(0.010222655652, 0.000818485952),
    to_complex(0.002286752946, - 0.014754814636),
    to_complex(0.001060069591, - 0.001662133807),
    to_complex(0.005933455360, - 0.006840245924),
    to_complex(0.002197903363, 0.001124132291),
    to_complex(0.000411028190, 0.007393274698),
    to_complex(0.014363410450, 0.002016585538),
    to_complex(0.005146056862, - 0.015672793855),
    to_complex(0.008623650342, - 0.007989113731),
    to_complex(0.000895303135, - 0.018844312607),
    to_complex(0.012676689064, - 0.003792693192),
    to_complex(- 0.016652906889, - 0.012520422771),
    to_complex(0.007079997943, - 0.002509704072),
    to_complex(- 0.003868765883, - 0.005401615113),
    to_complex(- 0.006873706323, - 0.005311525982),
    to_complex(- 0.009603924149, 0.005366157679),
    to_complex(0.004984735012, 0.012541472827),
    to_complex(- 0.001792377047, 0.014580420749),
    to_complex(- 0.003142233997, 0.015046392583),
    to_complex(0.003092203234, - 0.008940502572),
    to_complex(0.002620038037, - 0.000734151772),
    to_complex(- 0.000928615698, 0.017657556983),
    to_complex(0.006733799209, 0.002656892281),
    to_complex(- 0.007756596641, - 0.015750473767),
    to_complex(0.009182601659, 0.001333416849),
    to_complex(- 0.003535236039, - 0.004299879651),
    to_complex(- 0.001596831507, 0.012134040221),
    to_complex(0.003696910498, 0.009285595914),
    to_complex(0.008524870081, 0.004907594512),
    to_complex(0.001839513859, - 0.007734644188),
    to_complex(0.003877413966, 0.007385696685),
    to_complex(0.004057370040, 0.003228870754),
    to_complex(0.013002438135, - 0.003121934768),
    to_complex(- 0.002447720621, - 0.003258238945),
    to_complex(0.004552170841, 0.006054753457),
    to_complex(0.012249806442, - 0.010695602138),
    to_complex(0.001174520739, - 0.010008800858),
    to_complex(0.000680446592, - 0.007145296853),
    to_complex(0.003104168375, - 0.002072261105),
    to_complex(0.013686862742, 0.001925796801),
    to_complex(- 0.002325916830, - 0.013015627111),
    to_complex(0.009283385981, 0.001592941565),
    to_complex(0.001390659010, - 0.008899421081),
    to_complex(- 0.004431196053, 0.002408969961),
    to_complex(0.001076077423, 0.002799488578),
    to_complex(- 0.004594026817, 0.003146228111),
    to_complex(- 0.008325207132, 0.006612510465),
    to_complex(- 0.002018742091, - 0.001337435618),
    to_complex(0.001775452607, - 0.006134194178),
    to_complex(0.010978951834, 0.005931461915),
    to_complex(0.008432310972, 0.010410314306),
    to_complex(0.000315297868, - 0.005364185056),
    to_complex(0.008021507185, - 0.010193063925),
    to_complex(0.002906680338, - 0.001794823417),
    to_complex(0.007522908566, 0.017890432960),
    to_complex(0.006121369481, - 0.003887830885),
    to_complex(- 0.012353390582, - 0.006058673838),
    to_complex(- 0.009604983923, - 0.003164207565),
    to_complex(- 0.003692809107, - 0.005526282792),
    to_complex(0.006582459965, - 0.008618183552),
    to_complex(0.014016487821, 0.003701457743),
    to_complex(- 0.005567779464, 0.007169589798),
    to_complex(0.002343207034, - 0.008902211410),
    to_complex(- 0.001794298942, - 0.009414403283),
    to_complex(0.009234078328, 0.011344128503),
    to_complex(0.008394552721, 0.007734999526),
    to_complex(- 0.003044973324, - 0.001324633083),
    to_complex(0.014698265718, - 0.007741348127),
    to_complex(0.003010240727, - 0.000103380214),
    to_complex(- 0.003615131911, 0.003666638355),
    to_complex(0.005348611687, 0.004327837456),
    to_complex(- 0.003571929591, - 0.010714841127),
    to_complex(- 0.000975695761, 0.011559489815),
    to_complex(- 0.004044050388, - 0.002710609933),
    to_complex(0.008305945440, 0.010735421262),
    to_complex(- 0.000502030209, 0.002161492100),
    to_complex(0.005121564099, 0.001066662641),
    to_complex(0.003949640732, - 0.000921512515),
    to_complex(- 0.004746149567, - 0.004263943396),
    to_complex(0.010904017201, - 0.015302768076),
    to_complex(0.000849287733, - 0.007495860455),
    to_complex(0.009250865105, 0.007766647889),
    to_complex(0.009694179420, 0.008543159870),
    to_complex(- 0.016669076830, - 0.002088961554),
    to_complex(0.002594047692, - 0.003076499876),
    to_complex(0.000466693988, 0.005182497940),
    to_complex(0.010176487035, 0.006414408495),
    to_complex(0.002998029209, - 0.011472975166),
    to_complex(0.007876820465, 0.006954795614),
    to_complex(- 0.007854676940, 0.002651117629),
    to_complex(0.001720015383, 0.000246334117),
    to_complex(0.005335365743, - 0.001304569509),
    to_complex(0.019403163614, - 0.001125933817),
    to_complex(- 0.004047900475, 0.000252173838),
    to_complex(- 0.004012593163, 0.005875268194),
    to_complex(0.004742927309, 0.000525593937),
    to_complex(0.002107865769, 0.009410434009),
    to_complex(0.004139173598, 0.002650256293),
    to_complex(0.000798724739, - 0.009863283123),
    to_complex(- 0.006732760861, 0.002574148969),
    to_complex(0.006032655079, - 0.003023837708),
    to_complex(0.002608517657, - 0.006702558019),
    to_complex(- 0.005309076535, - 0.002625169867),
    to_complex(- 0.000167943903, 0.006063012205),
    to_complex(- 0.004280948030, - 0.008668212544),
    to_complex(- 0.002014441559, 0.006054479710),
    to_complex(- 0.009594365216, - 0.002887562818),
    to_complex(0.005362076894, - 0.004278177703),
    to_complex(0.005637001526, - 0.004921125760),
    to_complex(0.008925021507, - 0.001071228187),
    to_complex(- 0.006216298587, 0.007640954981),
    to_complex(0.012085288538, - 0.004561026738),
    to_complex(0.004625649356, - 0.000179514503),
    to_complex(- 0.005450114969, - 0.007053517272),
    to_complex(- 0.005294967787, - 0.007299741368),
    to_complex(- 0.004814398472, - 0.003305479816),
    to_complex(0.006178589423, 0.004189210226),
    to_complex(- 0.001024223868, 0.002084577196),
    to_complex(- 0.015872508668, - 0.004878460637),
    to_complex(- 0.003219743001, - 0.003336181353),
    to_complex(0.004636112095, 0.006692967921),
    to_complex(0.012141503757, 0.000316308433),
    to_complex(0.005228368622, 0.010546483130),
    to_complex(- 0.005825574894, - 0.008214421643),
    to_complex(0.002539752390, - 0.009674765002),
    to_complex(0.017002335029, 0.003829914882),
    to_complex(0.006511965032, - 0.002844918109),
    to_complex(0.006990817118, - 0.002456147423),
    to_complex(0.012903098309, 0.001213705470),
    to_complex(- 0.007866412794, 0.013099136816),
    to_complex(- 0.005469299667, - 0.007505318705),
    to_complex(0.000267218008, 0.000006492430),
    to_complex(0.013622442975, 0.007768623124),
    to_complex(- 0.003986811010, - 0.003573432190),
    to_complex(- 0.000582697840, - 0.000283488478),
    to_complex(0.003246418584, 0.006610687301),
    to_complex(0.017243259127, - 0.006568966786),
    to_complex(0.008939994202, 0.004507149270),
    to_complex(- 0.003725267381, - 0.003192691042),
    to_complex(- 0.001180786198, 0.000250669703),
    to_complex(0.002569702867, 0.005478109419),
    to_complex(- 0.004228165308, 0.016167928026),
    to_complex(- 0.002039615891, - 0.010969039525),
    to_complex(- 0.003674510616, - 0.000178512008),
    to_complex(0.000452234258, - 0.001282633007),
    to_complex(- 0.001623311047, - 0.000112917141),
    to_complex(- 0.009201396506, - 0.002744818451),
    to_complex(0.006425573898, - 0.011017677109),
    to_complex(0.006630303148, 0.000381782378),
    to_complex(- 0.003459623800, 0.005593643672),
    to_complex(0.012659048394, - 0.001195491878),
    to_complex(- 0.002481692524, 0.016340553588),
    to_complex(0.013680194081, - 0.011260458084),
    to_complex(- 0.002997757876, 0.002507658155),
    to_complex(- 0.003789797728, 0.010280353826),
    to_complex(- 0.007377153378, - 0.010824617659),
    to_complex(0.016871577772, - 0.010863992549),
    to_complex(- 0.000771234905, 0.002883632203),
    to_complex(- 0.014700995713, - 0.004492714053),
    to_complex(0.006120397404, - 0.007405663385),
    to_complex(0.005067373496, - 0.009101667254),
    to_complex(0.012405596061, 0.005513062403),
    to_complex(0.008640597394, - 0.010125186008),
    to_complex(- 0.013362727373, - 0.003188958913),
    to_complex(0.013411339016, - 0.010124257739),
    to_complex(0.009599661895, 0.001055060656),
    to_complex(- 0.008986306000, - 0.006616504583),
    to_complex(0.009816568508, 0.006791814416),
    to_complex(0.006455058949, - 0.000854448909),
    to_complex(0.009735066801, 0.008386096877),
    to_complex(0.000794233158, - 0.006093245972),
    to_complex(- 0.008305551020, 0.003414034856),
    to_complex(0.011914903984, 0.012365849089),
    to_complex(0.002081818846, - 0.012047437785),
    to_complex(- 0.003455714977, - 0.002369015706),
    to_complex(- 0.002022972490, - 0.001600927876),
    to_complex(- 0.000239432680, - 0.007660896388),
    to_complex(0.004039397559, 0.016754580470),
    to_complex(0.011246502874, - 0.001118547370),
    to_complex(- 0.006379097687, 0.011090121954),
    to_complex(0.012231057268, - 0.007100165708),
    to_complex(- 0.000491341425, 0.000301779707),
    to_complex(- 0.005022674841, - 0.003775297130),
    to_complex(0.002294618827, - 0.018908959185),
    to_complex(0.000818537791, - 0.005758286140),
    to_complex(- 0.005500775665, - 0.000932140016),
    to_complex(- 0.001918094188, 0.000643959906),
    to_complex(- 0.009962721320, - 0.012946350632),
    to_complex(0.008201928159, 0.000534217581),
    to_complex(0.000475569825, 0.006698527808),
    to_complex(0.008977850450, 0.002356138966),
    to_complex(0.013255258459, - 0.001926500573),
    to_complex(0.015613200014, 0.002557172398),
    to_complex(- 0.000049170732, 0.006218671265),
    to_complex(0.001144114771, - 0.003014032837),
    to_complex(0.004791457089, - 0.000668932223),
    to_complex(0.008927797265, 0.007998612910),
    to_complex(0.002330716898, - 0.007605195510),
    to_complex(- 0.004885160873, 0.006826892157),
    to_complex(- 0.003247705305, 0.000757886735),
    to_complex(0.016419710546, 0.013349598739),
    to_complex(0.002069052381, 0.005637627210),
    to_complex(- 0.004691591883, 0.002714949811),
    to_complex(0.002573797190, - 0.006277565429),
    to_complex(0.010492620169, 0.012447067454),
    to_complex(0.004516306745, - 0.002358650343),
    to_complex(0.001196752444, - 0.004314753409),
    to_complex(- 0.007372709740, - 0.004173719236),
    to_complex(- 0.003256459409, - 0.000124791524),
    to_complex(0.008274175372, - 0.005715765499),
    to_complex(0.000659257880, 0.001025635700),
    to_complex(- 0.010053369658, - 0.004733410330),
    to_complex(0.005576561314, 0.012028694649),
    to_complex(- 0.009277843627, - 0.000575228342),
    to_complex(0.004976927472, - 0.002386627457),
    to_complex(0.008908612854, 0.005980466854),
    to_complex(0.003198639904, - 0.003178178762),
    to_complex(0.001104432377, 0.007893369337),
    to_complex(0.009152076606, 0.000158229664),
    to_complex(0.004590110289, - 0.011489743987),
    to_complex(0.008626385347, - 0.004091824372),
    to_complex(- 0.001445056260, 0.001905576269),
    to_complex(0.003903959328, 0.003081041142),
    to_complex(- 0.000967407543, 0.011185563355),
    to_complex(0.011533488712, 0.001346675955),
    to_complex(- 0.004176667424, 0.009106353585),
    to_complex(- 0.001228532582, - 0.005888464228),
    to_complex(0.008351271805, - 0.009285130337),
    to_complex(- 0.002996429740, - 0.004590702064),
    to_complex(0.004068481671, 0.002868069018),
    to_complex(- 0.006330802954, 0.002205354201),
    to_complex(0.001370612936, - 0.010333705923),
    to_complex(0.007195813499, - 0.004465856805),
    to_complex(0.008576066093, 0.017727496016),
    to_complex(- 0.000994610117, 0.003814499872),
    to_complex(0.005528766161, 0.004289025192),
    to_complex(0.000145202146, - 0.010309205297),
    to_complex(- 0.001935066694, 0.001639690536),
    to_complex(- 0.004803521338, - 0.011030233995),
    to_complex(0.000409938656, - 0.002740425071),
    to_complex(0.007051870563, 0.000450488983),
    to_complex(- 0.010392005159, 0.012319602574),
    to_complex(- 0.004558163847, - 0.002135736414),
    to_complex(0.003778847712, 0.003871847346),
    to_complex(0.005596377018, - 0.007192939791),
    to_complex(0.008106474005, - 0.008354078295),
    to_complex(- 0.006742923336, 0.009511377763),
    to_complex(0.005020665513, 0.001697154856),
    to_complex(0.002734721179, 0.005832783124),
    to_complex(0.002735791722, 0.004360039810),
    to_complex(- 0.006119901805, - 0.010503949312),
    to_complex(- 0.001150240843, 0.002426581065),
    to_complex(0.014294911916, - 0.000957821453),
    to_complex(- 0.002420041353, 0.003925982225),
    to_complex(- 0.003238642165, 0.000777485406),
    to_complex(0.005955032834, - 0.010427584085),
    to_complex(0.014246515155, 0.004566647614),
    to_complex(0.000816066920, - 0.002421778079),
    to_complex(- 0.008594930710, - 0.000872754068),
    to_complex(- 0.003029344458, - 0.010429835124),
    to_complex(0.010556577542, - 0.006656808579),
    to_complex(0.011517057169, - 0.016013681994),
    to_complex(- 0.015211476518, 0.003048172104),
    to_complex(0.007770822174, - 0.004435631387),
    to_complex(0.013373596257, 0.001720597622),
    to_complex(0.012540141897, - 0.005581448860),
    to_complex(0.003898078330, - 0.003766014236),
    to_complex(- 0.002836827788, - 0.008962881754),
    to_complex(0.017539910921, - 0.005786903112),
    to_complex(- 0.000370711449, 0.001932416429),
    to_complex(- 0.006912097094, 0.001000344860),
    to_complex(0.007765164358, - 0.000973142528),
    to_complex(0.010164772900, 0.009230222065),
    to_complex(- 0.001530823338, 0.010344035742),
    to_complex(- 0.001595738391, 0.000165253631),
    to_complex(- 0.006625528841, - 0.002254661542),
    to_complex(0.017412267750, 0.000579061437),
    to_complex(- 0.011787897886, 0.003527961834),
    to_complex(0.004941665914, 0.007004421941),
    to_complex(0.003534235741, 0.007375657127),
    to_complex(0.011280011057, 0.000935413647),
    to_complex(0.005349576400, 0.006634579079),
    to_complex(- 0.012364229325, - 0.001509633787),
    to_complex(0.004898114038, - 0.017328486000),
    to_complex(0.005620209675, - 0.000813002004),
    to_complex(0.005803146590, - 0.011555070895),
    to_complex(- 0.016812401483, - 0.003194330036),
    to_complex(0.003478290054, 0.011969850456),
    to_complex(- 0.005773131419, 0.006050798137),
    to_complex(- 0.001739675826, - 0.006947083155),
    to_complex(0.006028172365, - 0.003059060094),
    to_complex(0.004913735427, - 0.003444707901),
    to_complex(0.006217043748, - 0.009497303643),
    to_complex(0.004818796594, 0.002689738170),
    to_complex(- 0.004479695655, 0.001392524871),
    to_complex(- 0.001367643862, - 0.006796381618),
    to_complex(0.013086067744, - 0.004223003753),
    to_complex(0.005029691374, 0.005745173498),
    to_complex(- 0.004642755149, 0.004864622872),
    to_complex(- 0.002060879935, - 0.001842057289),
    to_complex(- 0.002316530112, - 0.004602486827),
    to_complex(- 0.000529281862, 0.008560576504),
    to_complex(- 0.002016293287, - 0.001525788338),
    to_complex(0.009352053405, - 0.001855991777),
    to_complex(0.010664489743, 0.002631819773),
    to_complex(0.004029329335, 0.006536894055),
    to_complex(0.000497245737, 0.005118258465),
    to_complex(0.001082982132, - 0.004368546324),
    to_complex(0.005624460000, 0.010120922732),
    to_complex(0.003877319905, 0.002025348043),
    to_complex(- 0.002823672470, - 0.000934240074),
    to_complex(0.001759497304, - 0.002807271349),
    to_complex(0.021246200454, - 0.009409115899),
    to_complex(0.004655002529, 0.000456970090),
    to_complex(0.003079708479, 0.003567851944),
    to_complex(- 0.005950314090, 0.004339535286),
    to_complex(0.019553315017, - 0.013164512719),
    to_complex(0.000124100066, 0.001615368168),
    to_complex(- 0.005690969062, - 0.009652772405),
    to_complex(- 0.005373524378, - 0.019028034326),
    to_complex(0.017427945074, 0.007005601155),
    to_complex(0.007736744504, 0.009301620182),
    to_complex(0.007822400992, - 0.000830520450),
    to_complex(- 0.006988740410, 0.010018082757),
    to_complex(0.005198075771, - 0.002426556992),
    to_complex(- 0.001488003750, 0.006058090829),
    to_complex(- 0.005333030450, 0.004119934597),
    to_complex(- 0.004239908245, - 0.005377636931),
    to_complex(0.004431355481, - 0.014690046778),
    to_complex(- 0.003284564642, 0.007016580948),
    to_complex(0.000781227006, - 0.000506051543),
    to_complex(0.000665615153, - 0.011922887872),
    to_complex(- 0.002790354355, - 0.007095106460),
    to_complex(0.000298008590, 0.005107250417),
    to_complex(- 0.004687856475, - 0.008448301707),
    to_complex(0.000096804435, - 0.008226159217),
    to_complex(0.016697290188, - 0.001417636768),
    to_complex(0.003242876098, 0.004068573483),
    to_complex(- 0.010054936536, - 0.004857048982),
    to_complex(- 0.004810612030, - 0.003657769865),
    to_complex(- 0.001493545652, 0.001633319216),
    to_complex(0.000487115935, - 0.006899753766),
    to_complex(- 0.007334422232, 0.001401612163),
    to_complex(0.000154717718, - 0.001322627957),
    to_complex(0.006005603876, - 0.007120846565),
    to_complex(- 0.001341682203, 0.000061064644),
    to_complex(- 0.009138750223, - 0.002057491521),
    to_complex(- 0.003496249805, - 0.004635437643),
    to_complex(0.006526293733, - 0.007199299992),
    to_complex(0.008925460010, 0.005967666900),
    to_complex(0.004787419484, 0.004814971464),
    to_complex(0.007506481952, - 0.008480506143),
    to_complex(0.016152021368, 0.001597014881),
    to_complex(0.009566912809, - 0.008448053348),
    to_complex(- 0.002575675187, - 0.001702976171),
    to_complex(- 0.007795400047, - 0.000472931598),
    to_complex(0.020441114217, - 0.010698053261),
    to_complex(- 0.003712193101, 0.009583406349),
    to_complex(0.006445149610, - 0.004749603268),
    to_complex(0.001702053893, - 0.012548769541),
    to_complex(0.015292795931, 0.007431116307),
    to_complex(0.010194677701, 0.007370338225),
    to_complex(- 0.004539427823, 0.006333954614),
    to_complex(- 0.012298163044, 0.022788344898),
    to_complex(0.014336584522, - 0.013955229554),
    to_complex(- 0.006326594378, 0.007351425858),
    to_complex(- 0.012343128272, 0.000247685636),
    to_complex(- 0.002377827008, 0.006250976027),
    to_complex(0.022124005650, 0.006332616786),
    to_complex(- 0.008220290199, 0.011704480891),
    to_complex(- 0.001105555319, 0.002664337533),
    to_complex(- 0.000784686632, - 0.011165467267),
    to_complex(0.002548366920, - 0.009253482532),
    to_complex(0.004711461272, 0.005551381886),
    to_complex(- 0.010403868888, 0.007248580867),
    to_complex(0.004901836174, 0.009808380043),
    to_complex(0.006907973327, - 0.018573514421),
    to_complex(- 0.005409265023, - 0.005228234363),
    to_complex(- 0.005907005227, - 0.000779828207),
    to_complex(0.002800986892, 0.007095911222),
    to_complex(0.010913776828, - 0.011098809717),
    to_complex(0.007954259275, 0.008665577479),
    to_complex(- 0.002968338562, - 0.000912171715),
    to_complex(- 0.000115068172, 0.009967208255),
    to_complex(0.004438676158, - 0.000238693804),
    to_complex(0.022695097025, 0.000578080811),
    to_complex(0.009807994469, - 0.001282473214),
    to_complex(0.000145416808, 0.003596541587),
    to_complex(0.011478162008, 0.002575868361),
    to_complex(0.005823480400, 0.004941892272),
    to_complex(0.003336274678, 0.012544919408),
    to_complex(- 0.005526148214, - 0.007209206120),
    to_complex(- 0.001981738865, 0.009896727535),
    to_complex(0.005929906801, - 0.003057078985),
    to_complex(- 0.005546519307, - 0.003034588487),
    to_complex(0.005576576638, 0.007967615750),
    to_complex(0.023449215040, - 0.004186941115),
    to_complex(- 0.005767832761, - 0.000653029940),
    to_complex(0.007123200170, 0.001326836551),
    to_complex(0.002582199735, - 0.008045729083),
    to_complex(0.018242245637, 0.003433652436),
    to_complex(0.005314745031, - 0.004312318827),
    to_complex(0.012636494097, - 0.008368640563),
    to_complex(- 0.001679492666, - 0.002383731244),
    to_complex(0.019151624031, - 0.001661308164),
    to_complex(0.004871650292, 0.002734864486),
    to_complex(- 0.015711638471, 0.001997280222),
    to_complex(- 0.009250011290, - 0.006800660769),
    to_complex(0.005545511569, - 0.003317621794),
    to_complex(0.009320581690, - 0.001777780243),
    to_complex(0.001353830474, 0.017015400703),
    to_complex(- 0.014041165867, - 0.004884122984),
    to_complex(0.011177249312, - 0.010367923795),
    to_complex(- 0.000982965345, 0.005173276534),
    to_complex(- 0.001166721873, 0.004361251904),
    to_complex(0.004012323022, 0.003834820594),
    to_complex(0.005318245866, - 0.001358031159),
    to_complex(- 0.001185596702, 0.018504250136),
    to_complex(0.011278237377, - 0.002170327420),
    to_complex(- 0.002898694300, 0.010797416049),
    to_complex(0.028641241507, 0.004383184044),
    to_complex(- 0.001847033074, 0.008836220181),
    to_complex(0.005036052392, - 0.005977957123),
    to_complex(0.000655947815, - 0.006599470654),
    to_complex(0.007634618164, - 0.005020684617),
    to_complex(- 0.004528714198, 0.009795886434),
    to_complex(0.008627144478, 0.001307402037),
    to_complex(- 0.007851386842, 0.000032972150),
    to_complex(0.011010455064, - 0.008114547083),
    to_complex(- 0.007314147750, 0.005160226240),
    to_complex(0.006121440419, - 0.006254081384),
    to_complex(0.006712625405, - 0.005866625460),
    to_complex(0.006575117872, 0.003572983824),
    to_complex(0.017695338175, 0.006701602652),
    to_complex(- 0.002005498655, - 0.013139452216),
    to_complex(- 0.003026171148, 0.000684132677),
    to_complex(0.021113461557, - 0.009868982303),
    to_complex(- 0.010445329626, 0.002425784300),
    to_complex(0.001608814165, 0.009468239828),
    to_complex(0.003346426717, 0.004875826845),
    to_complex(0.015307043206, - 0.013762245286),
    to_complex(0.004210630015, 0.011986321661),
    to_complex(0.005273882437, - 0.017753157434),
    to_complex(- 0.003148178229, - 0.001696080809),
    to_complex(0.014125834923, - 0.002055121277),
    to_complex(- 0.007548015196, - 0.006998892746),
    to_complex(0.001590631223, 0.012540849316),
    to_complex(0.000507570216, - 0.000031822525),
    to_complex(0.020861153811, - 0.016322793266),
    to_complex(0.006780683359, - 0.006783485639),
    to_complex(- 0.006134172395, - 0.002154919922),
    to_complex(0.002043737439, 0.009923172331),
    to_complex(0.023016082654, - 0.006311449842),
    to_complex(- 0.004877593876, - 0.003119817103),
    to_complex(0.006555681563, - 0.007741975624),
    to_complex(0.010376576815, - 0.010677030314),
    to_complex(0.011817921786, - 0.012322610562),
    to_complex(0.005333657663, 0.009950080644),
    to_complex(0.001060166409, 0.003618462894),
    to_complex(- 0.005132024760, - 0.010087689967),
    to_complex(0.012466373742, - 0.010720690546),
    to_complex(- 0.002662075421, 0.006623285938),
    to_complex(- 0.010059618337, - 0.001046152874),
    to_complex(- 0.008059405559, - 0.013072658773),
    to_complex(0.003722645810, - 0.009062482809),
    to_complex(0.005230782345, 0.002265232967),
    to_complex(0.010298613989, - 0.000075170492),
    to_complex(- 0.004472440144, 0.004088455950),
    to_complex(0.010304262033, 0.008808905016),
    to_complex(0.004554064004, 0.009465642245),
    to_complex(0.002092651825, 0.005191360045),
    to_complex(- 0.008298896314, 0.003688269515),
    to_complex(0.013549220058, - 0.017571879943),
    to_complex(0.007526279960, 0.010034135637),
    to_complex(0.006067419563, - 0.001773746331),
    to_complex(0.001684779245, - 0.002744298681),
    to_complex(0.011437888787, - 0.018802180052),
    to_complex(- 0.005779114854, 0.015448300295),
    to_complex(0.000657618128, - 0.000268660219),
    to_complex(0.001477503004, - 0.006676609736),
    to_complex(0.012837711465, - 0.007606743853),
    to_complex(0.010691551803, 0.011815859982),
    to_complex(0.005446173340, 0.005508444265),
    to_complex(- 0.002985617851, 0.004344778531),
    to_complex(0.019437505190, 0.000084167710),
    to_complex(0.004665255907, 0.005397607679),
    to_complex(- 0.006597113133, - 0.001182403336),
    to_complex(- 0.009629345968, 0.002296122733),
    to_complex(0.026387759889, - 0.010853424384),
    to_complex(0.004512348010, 0.001746367719),
    to_complex(0.000531629007, 0.005072332415),
    to_complex(- 0.004435887620, 0.000332198880),
    to_complex(0.008827061699, - 0.006195885754),
    to_complex(0.005913001809, 0.002293281192),
    to_complex(- 0.001925767264, - 0.005236607979),
    to_complex(- 0.008904628618, - 0.005441559131),
    to_complex(0.030186905381, - 0.003620144277),
    to_complex(0.004247330211, - 0.015065654208),
    to_complex(0.002465839164, - 0.010965170533),
    to_complex(- 0.008523595156, 0.005029475791),
    to_complex(0.021431895352, - 0.012512664924),
    to_complex(0.001463122118, - 0.001042234978),
    to_complex(0.002368774715, 0.007271767642),
    to_complex(0.001663302261, - 0.015294060227),
    to_complex(0.027865903183, - 0.014843006590),
    to_complex(- 0.005387327049, 0.006022316285),
    to_complex(- 0.007414061849, - 0.003683880991),
    to_complex(0.004457057973, - 0.001742795049),
    to_complex(0.021956837796, - 0.006768769984),
    to_complex(- 0.000581994344, 0.000632201811),
    to_complex(- 0.002050346880, - 0.014881422192),
    to_complex(0.002068677056, - 0.008564682783),
    to_complex(0.017229937229, - 0.022755747802),
    to_complex(0.014330280024, - 0.000556246747),
    to_complex(0.004677543424, - 0.009336132347),
    to_complex(- 0.015144212688, - 0.003901748575),
    to_complex(0.016991072061, - 0.007378745156),
    to_complex(0.000589790098, 0.003458122323),
    to_complex(0.007630737413, - 0.000250331890),
    to_complex(- 0.002091465440, 0.000503798031),
    to_complex(0.009016682113, - 0.015491343992),
    to_complex(0.001647357983, 0.012801461882),
    to_complex(0.010979951685, - 0.003137016118),
    to_complex(- 0.004038410356, - 0.001911611355),
    to_complex(0.012859899782, - 0.012089958198),
    to_complex(0.005291854769, 0.000502630258),
    to_complex(0.011716390282, - 0.000599429568),
    to_complex(- 0.000799325327, - 0.001631086182),
    to_complex(0.010959792409, - 0.014816322542),
    to_complex(0.009912772637, - 0.002695036705),
    to_complex(0.014814496598, 0.000511852126),
    to_complex(0.002675874354, - 0.005628676393),
    to_complex(0.027706603203, - 0.015942304188),
    to_complex(- 0.000904213510, - 0.000952461753),
    to_complex(- 0.004139637485, 0.000113489781),
    to_complex(- 0.009764242039, - 0.001570257746),
    to_complex(0.016937931778, 0.007116364990),
    to_complex(- 0.001345827612, 0.012884143175),
    to_complex(0.005896214424, 0.015206818229),
    to_complex(- 0.004073433760, - 0.006746279317),
    to_complex(0.028816309305, - 0.011980123552),
    to_complex(0.005563771759, 0.009251364794),
    to_complex(- 0.000034985934, - 0.005783922766),
    to_complex(- 0.014807449035, - 0.014452854805),
    to_complex(0.014497123347, - 0.023582465744),
    to_complex(0.009957646882, - 0.003482814383),
    to_complex(0.001526823231, - 0.003487046676),
    to_complex(- 0.003396082218, - 0.009464310852),
    to_complex(0.024195906577, - 0.010201550914),
    to_complex(- 0.003164840802, 0.004740286184),
    to_complex(0.000014788323, - 0.008524411815),
    to_complex(- 0.008474012195, - 0.015298019993),
    to_complex(0.017497476584, - 0.012330596533),
    to_complex(0.008405431215, - 0.005121338673),
    to_complex(0.007394357187, - 0.000047068287),
    to_complex(0.001425433874, 0.000800280639),
    to_complex(0.033310809233, - 0.021721551999),
    to_complex(0.003614899063, 0.013061152637),
    to_complex(- 0.005569496091, 0.003460439526),
    to_complex(- 0.004293446466, - 0.009246381658),
    to_complex(0.019205757239, - 0.018650103380),
    to_complex(0.000763020917, 0.014349891109),
    to_complex(0.001835421023, - 0.002248125723),
    to_complex(- 0.005626806483, - 0.018720311774),
    to_complex(0.036606395710, - 0.031348492597),
    to_complex(- 0.001623121635, 0.009773235077),
    to_complex(0.003198314753, 0.000852772802),
    to_complex(- 0.007336070659, - 0.011753761148),
    to_complex(0.021137051010, - 0.019343316838),
    to_complex(0.002155938292, 0.004631905182),
    to_complex(0.002581368203, 0.006375822851),
    to_complex(- 0.016802867993, 0.001195612915),
    to_complex(0.026640990919, - 0.019023289361),
    to_complex(- 0.000123136528, - 0.000254215045),
    to_complex(- 0.003741244536, 0.001360876505),
    to_complex(0.002121625160, 0.004746311460),
    to_complex(0.038663028779, - 0.019012181812),
    to_complex(- 0.007190577163, 0.005932501172),
    to_complex(- 0.004221350811, - 0.000762310291),
    to_complex(- 0.003708797083, - 0.016539685627),
    to_complex(0.028308543354, - 0.019690040002),
    to_complex(0.009527345765, 0.009370334165),
    to_complex(0.000794889798, - 0.020744510215),
    to_complex(- 0.011476614215, - 0.018656840579),
    to_complex(0.030731497343, - 0.018618471432),
    to_complex(- 0.003656349139, 0.005909295916),
    to_complex(- 0.003285500845, - 0.001424345423),
    to_complex(0.002294222179, - 0.006851179797),
    to_complex(0.026490672626, - 0.030105831521),
    to_complex(0.012769006712, 0.008149095307),
    to_complex(0.005166527275, 0.005267590226),
    to_complex(- 0.004027190142, - 0.016211553466),
    to_complex(0.036026934442, - 0.020305407629),
    to_complex(0.007049014584, 0.003023996984),
    to_complex(0.004723216372, 0.004389889471),
    to_complex(- 0.001558781326, - 0.003040610658),
    to_complex(0.022574137916, - 0.015479476225),
    to_complex(0.009873086148, 0.012633701220),
    to_complex(- 0.008944049662, - 0.001431941447),
    to_complex(- 0.002228757063, - 0.004053629769),
    to_complex(0.040307986154, - 0.022798217618),
    to_complex(0.005449313443, 0.007814338232),
    to_complex(- 0.007994176579, 0.006435096054),
    to_complex(- 0.017618952767, - 0.001785826893),
    to_complex(0.039928807907, - 0.033342689400),
    to_complex(- 0.005545175620, 0.010223276563),
    to_complex(0.001743292285, 0.000014482194),
    to_complex(- 0.010876499487, 0.003048564431),
    to_complex(0.035168355082, - 0.036433377087),
    to_complex(0.004356902223, 0.005181162200),
    to_complex(- 0.001782196234, - 0.013327838629),
    to_complex(0.004141734696, - 0.021873532882),
    to_complex(0.044444181603, - 0.013826733956),
    to_complex(0.015004230583, 0.010624693422),
    to_complex(0.005680260354, 0.009586948900),
    to_complex(- 0.009298717920, - 0.013779450150),
    to_complex(0.033979170596, - 0.031965688450),
    to_complex(0.011838259417, 0.001750919236),
    to_complex(- 0.017054585138, - 0.016004032744),
    to_complex(0.003045510935, 0.003825175874),
    to_complex(0.044371930109, - 0.033642538160),
    to_complex(0.014678064263, 0.005254658884),
    to_complex(0.004010000314, - 0.000537918292),
    to_complex(- 0.012074013593, 0.001074222258),
    to_complex(0.032551990358, - 0.036357652409),
    to_complex(0.014455725822, 0.023168621477),
    to_complex(- 0.011390643749, - 0.001584084973),
    to_complex(- 0.014897356748, - 0.017286270415),
    to_complex(0.048939291238, - 0.029474702568),
    to_complex(0.009268415809, - 0.002047289446),
    to_complex(- 0.000444148577, 0.005817010398),
    to_complex(0.002509924074, - 0.002315797175),
    to_complex(0.048139689361, - 0.043604827418),
    to_complex(0.018300822184, 0.018753170714),
    to_complex(0.002802829885, 0.012863223213),
    to_complex(- 0.004262746820, - 0.015219728872),
    to_complex(0.055522722166, - 0.046242068531),
    to_complex(0.003591235495, 0.014540980968),
    to_complex(- 0.002784254556, - 0.004077659569),
    to_complex(- 0.009984947863, 0.002997739358),
    to_complex(0.057922010029, - 0.052448353016),
    to_complex(0.010393287010, 0.025473594904),
    to_complex(- 0.020983473636, - 0.000426634948),
    to_complex(- 0.008483911314, - 0.016906264577),
    to_complex(0.061714171221, - 0.054078495913),
    to_complex(0.018244804257, 0.021070628679),
    to_complex(0.003468470115, - 0.006772633602),
    to_complex(- 0.012387720631, - 0.009359360318),
    to_complex(0.079227158055, - 0.058913055564),
    to_complex(0.023925350552, 0.017274972311),
    to_complex(0.005704025736, 0.004624671356),
    to_complex(- 0.031880490146, - 0.022111509628),
    to_complex(0.073851744519, - 0.065838505465),
    to_complex(0.024411241745, 0.008876664565),
    to_complex(0.002506405057, 0.001338020893),
    to_complex(- 0.024640828912, - 0.020370350345),
    to_complex(0.092572956150, - 0.076410575260),
    to_complex(0.022287391077, 0.033789596159),
    to_complex(- 0.004005816311, - 0.002607691371),
    to_complex(- 0.020227850693, - 0.017824641310),
    to_complex(0.098721974409, - 0.095633556706),
    to_complex(0.026974428989, 0.023851533795),
    to_complex(0.006203101104, - 0.002215837855),
    to_complex(- 0.027423747525, - 0.026790189785),
    to_complex(0.114007151945, - 0.122674393493),
    to_complex(0.043919100912, 0.028342759630),
    to_complex(- 0.004646280168, - 0.003295679855),
    to_complex(- 0.028458592098, - 0.048110001252),
    to_complex(0.146594493406, - 0.128814599440),
    to_complex(0.046864261896, 0.034286118288),
    to_complex(- 0.003182374439, - 0.003482134295),
    to_complex(- 0.041053397039, - 0.031124060265),
    to_complex(0.195468715643, - 0.175923894702),
    to_complex(0.045656287380, 0.047910872846),
    to_complex(- 0.006627592712, - 0.004121208884),
    to_complex(- 0.056271640358, - 0.047441938250),
    to_complex(0.260468640644, - 0.259310640181),
    to_complex(0.074157954230, 0.070121724177),
    to_complex(0.011433341872, 0.001002496238),
    to_complex(- 0.092355139255, - 0.097534905023),
    to_complex(0.419655691208, - 0.419001736817),
    to_complex(0.125889930241, 0.122552587264),
    to_complex(0.005885794485, 0.002408601835),
    to_complex(- 0.220700517194, - 0.213862796050),
    to_complex(1.274321145456, - 1.263756831848),
    to_complex(0.622618932598, 0.638254649110));

end input_data;
