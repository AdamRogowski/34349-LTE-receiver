library IEEE;
  use work.complex_pkg.all;

package input_data is

  constant INPUT_DATA_2048_16QAM_CLEAR : complex_array(0 to 2047) := (
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.637595835525, 0.635642710525),
    to_complex(- 1.269329299991, 1.277141799991),
    to_complex(- 0.213181655259, - 0.211228530259),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.128298020250, 0.126344895250),
    to_complex(- 0.420494947286, 0.428307447286),
    to_complex(- 0.091918748841, - 0.089965623841),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.071707598622, 0.069754473622),
    to_complex(- 0.250721684926, 0.258534184926),
    to_complex(- 0.058845594387, - 0.056892469387),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.049940822593, 0.047987697593),
    to_complex(- 0.177957149482, 0.185769649482),
    to_complex(- 0.043410390253, - 0.041457265253),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.038416295193, 0.036463170193),
    to_complex(- 0.137528856024, 0.145341356024),
    to_complex(- 0.034473378260, - 0.032520253260),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.031281302833, 0.029328177833),
    to_complex(- 0.111798854027, 0.119611354027),
    to_complex(- 0.028644197202, - 0.026691072202),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.026428868603, 0.024475743603),
    to_complex(- 0.093983316292, 0.101795816292),
    to_complex(- 0.024541588793, - 0.022588463793),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.022914485594, 0.020961360594),
    to_complex(- 0.080916456729, 0.088728956729),
    to_complex(- 0.021497202231, - 0.019544077231),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.020251589629, 0.018298464629),
    to_complex(- 0.070922270882, 0.078734770882),
    to_complex(- 0.019148218499, - 0.017195093499),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.018164022645, 0.016210897645),
    to_complex(- 0.063030440328, 0.070842940328),
    to_complex(- 0.017280667393, - 0.015327542393),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.016483395569, 0.014530270569),
    to_complex(- 0.056640291713, 0.064452791713),
    to_complex(- 0.015760195518, - 0.013807070518),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.015101190990, 0.013148065990),
    to_complex(- 0.051360081505, 0.059172581505),
    to_complex(- 0.014498186796, - 0.012545061796),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.013944325739, 0.011991200739),
    to_complex(- 0.046923424060, 0.054735924060),
    to_complex(- 0.013433826260, - 0.011480701260),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.012961779486, 0.011008654486),
    to_complex(- 0.043142862780, 0.050955362780),
    to_complex(- 0.012523990562, - 0.010570865562),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.012116853385, 0.010163728385),
    to_complex(- 0.039882653199, 0.047695153199),
    to_complex(- 0.011737250813, - 0.009784125813),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.011382474511, 0.009429349511),
    to_complex(- 0.037042081647, 0.044854581647),
    to_complex(- 0.011050160057, - 0.009097035057),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.010738234036, 0.008785109036),
    to_complex(- 0.034544849863, 0.042357349863),
    to_complex(- 0.010444870603, - 0.008491745603),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.010168455605, 0.008215330605),
    to_complex(- 0.032332099158, 0.040144599158),
    to_complex(- 0.009907556767, - 0.007954431767),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.009660898773, 0.007707773773),
    to_complex(- 0.030357697021, 0.038170197021),
    to_complex(- 0.009427342340, - 0.007474217340),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.009205866554, 0.007252741554),
    to_complex(- 0.028584973994, 0.036397473994),
    to_complex(- 0.008995553882, - 0.007042428882),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.008795577413, 0.006842452413),
    to_complex(- 0.026984415612, 0.034796915612),
    to_complex(- 0.008605189936, - 0.006652064936),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.008423714566, 0.006470589566),
    to_complex(- 0.025531998452, 0.033344498452),
    to_complex(- 0.008250536662, - 0.006297411662),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.008085096829, 0.006131971829),
    to_complex(- 0.024207969896, 0.032020469896),
    to_complex(- 0.007926884849, - 0.005973759849),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.007775434394, 0.005822309394),
    to_complex(- 0.022995939456, 0.030808439456),
    to_complex(- 0.007630318408, - 0.005677193408),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.007491145051, 0.005538020051),
    to_complex(- 0.021882192621, 0.029694692621),
    to_complex(- 0.007357554149, - 0.005404429149),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.007229214058, 0.005276089058),
    to_complex(- 0.020855166156, 0.028667666156),
    to_complex(- 0.007105818889, - 0.005152693889),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.006987086062, 0.005033961062),
    to_complex(- 0.019905042202, 0.027717542202),
    to_complex(- 0.006872754121, - 0.004919629121),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.006762580801, 0.004809455801),
    to_complex(- 0.019023430933, 0.026835930933),
    to_complex(- 0.006656341296, - 0.004703216296),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.006553826718, 0.004600701718),
    to_complex(- 0.018203120025, 0.026015620025),
    to_complex(- 0.006454842707, - 0.004501717707),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.006359208193, 0.004406083193),
    to_complex(- 0.017437875081, 0.025250375081),
    to_complex(- 0.006266754280, - 0.004313629280),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.006177323236, 0.004224198236),
    to_complex(- 0.016722279311, 0.024534779311),
    to_complex(- 0.006090767590, - 0.004137642590),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.006006949308, 0.004053824308),
    to_complex(- 0.016051603757, 0.023864103757),
    to_complex(- 0.005925739051, - 0.003972614051),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.005847015499, 0.003893890499),
    to_complex(- 0.015421701470, 0.023234201470),
    to_complex(- 0.005770664744, - 0.003817539744),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.005696579726, 0.003743454726),
    to_complex(- 0.014828920645, 0.022641420645),
    to_complex(- 0.005624659732, - 0.003671534732),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.005554809928, 0.003601684928),
    to_complex(- 0.014270032858, 0.022082532858),
    to_complex(- 0.005486940938, - 0.003533815938),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.005420968456, 0.003467843456),
    to_complex(- 0.013742173440, 0.021554673440),
    to_complex(- 0.005356812895, - 0.003403687895),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.005294399056, 0.003341274056),
    to_complex(- 0.013242791641, 0.021055291641),
    to_complex(- 0.005233655834, - 0.003280530834),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.005174515940, 0.003221390940),
    to_complex(- 0.012769608778, 0.020582108778),
    to_complex(- 0.005116915650, - 0.003163790650),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.005060794574, 0.003107669574),
    to_complex(- 0.012320582903, 0.020133082903),
    to_complex(- 0.005006095435, - 0.003052970435),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.004952763878, 0.002999638878),
    to_complex(- 0.011893878832, 0.019706378832),
    to_complex(- 0.004900748279, - 0.002947623279),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.004849999583, 0.002896874583),
    to_complex(- 0.011487842622, 0.019300342622),
    to_complex(- 0.004800471139, - 0.002847346139),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.004752118560, 0.002798993560),
    to_complex(- 0.011100979732, 0.018913479732),
    to_complex(- 0.004704899583, - 0.002751774583),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.004658773947, 0.002705648947),
    to_complex(- 0.010731936275, 0.018544436275),
    to_complex(- 0.004613703275, - 0.002660578275),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.004569650961, 0.002616525961),
    to_complex(- 0.010379482843, 0.018191982843),
    to_complex(- 0.004526582077, - 0.002573457077),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.004484463269, 0.002531338269),
    to_complex(- 0.010042500528, 0.017855000528),
    to_complex(- 0.004443262678, - 0.002490137678),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.004402949848, 0.002449824848),
    to_complex(- 0.009719968773, 0.017532468773),
    to_complex(- 0.004363495658, - 0.002410370658),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.004324872245, 0.002371747245),
    to_complex(- 0.009410954802, 0.017223454802),
    to_complex(- 0.004287052938, - 0.002333927938),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.004250012193, 0.002296887193),
    to_complex(- 0.009114604375, 0.016927104375),
    to_complex(- 0.004213725538, - 0.002260600538),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.004178169515, 0.002225044515),
    to_complex(- 0.008830133696, 0.016642633696),
    to_complex(- 0.004143321627, - 0.002190196627),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.004109160291, 0.002156035291),
    to_complex(- 0.008556822293, 0.016369322293),
    to_complex(- 0.004075664791, - 0.002122539791),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.004042815236, 0.002089690236),
    to_complex(- 0.008294006750, 0.016106506750),
    to_complex(- 0.004010592519, - 0.002057467519),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.003978978278, 0.002025853278),
    to_complex(- 0.008041075171, 0.015853575171),
    to_complex(- 0.003947954860, - 0.001994829860),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.003917505289, 0.001964380289),
    to_complex(- 0.007797462267, 0.015609962267),
    to_complex(- 0.003887613230, - 0.001934488230),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.003858262964, 0.001905137964),
    to_complex(- 0.007562645004, 0.015375145004),
    to_complex(- 0.003829439355, - 0.001876314355),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.003801127826, 0.001848002826),
    to_complex(- 0.007336138727, 0.015148638727),
    to_complex(- 0.003773314331, - 0.001820189331),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.003745985334, 0.001792860334),
    to_complex(- 0.007117493699, 0.014929993699),
    to_complex(- 0.003719127783, - 0.001766002783),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.003692729090, 0.001739604090),
    to_complex(- 0.006906292015, 0.014718792015),
    to_complex(- 0.003666777112, - 0.001713652112),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.003641260127, 0.001688135127),
    to_complex(- 0.006702144829, 0.014514644829),
    to_complex(- 0.003616166823, - 0.001663041823),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.003591486273, 0.001638361273),
    to_complex(- 0.006504689876, 0.014317189876),
    to_complex(- 0.003567207923, - 0.001614082923),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.003543321575, 0.001590196575),
    to_complex(- 0.006313589233, 0.014126089233),
    to_complex(- 0.003519817372, - 0.001566692372),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.003496685783, 0.001543560783),
    to_complex(- 0.006128527311, 0.013941027311),
    to_complex(- 0.003473917594, - 0.001520792594),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.003451503888, 0.001498378888),
    to_complex(- 0.005949209038, 0.013761709038),
    to_complex(- 0.003429436039, - 0.001476311039),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.003407705696, 0.001454580696),
    to_complex(- 0.005775358215, 0.013587858215),
    to_complex(- 0.003386304777, - 0.001433179777),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.003365225452, 0.001412100452),
    to_complex(- 0.005606716035, 0.013419216035),
    to_complex(- 0.003344460139, - 0.001391335139),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.003324001491, 0.001370876491),
    to_complex(- 0.005443039729, 0.013255539729),
    to_complex(- 0.003303842387, - 0.001350717387),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.003283975926, 0.001330850926),
    to_complex(- 0.005284101347, 0.013096601347),
    to_complex(- 0.003264395415, - 0.001311270415),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.003245094363, 0.001291969363),
    to_complex(- 0.005129686641, 0.012942186641),
    to_complex(- 0.003226066476, - 0.001272941476),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.003207305643, 0.001254180643),
    to_complex(- 0.004979594048, 0.012792094048),
    to_complex(- 0.003188805936, - 0.001235680936),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.003170561599, 0.001217436599),
    to_complex(- 0.004833633770, 0.012646133770),
    to_complex(- 0.003152567046, - 0.001199442046),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.003134816848, 0.001181691848),
    to_complex(- 0.004691626920, 0.012504126920),
    to_complex(- 0.003117305736, - 0.001164180736),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.003100028587, 0.001146903587),
    to_complex(- 0.004553404754, 0.012365904754),
    to_complex(- 0.003082980426, - 0.001129855426),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.003066156414, 0.001113031414),
    to_complex(- 0.004418807960, 0.012231307960),
    to_complex(- 0.003049551850, - 0.001096426850),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.003033162162, 0.001080037162),
    to_complex(- 0.004287686005, 0.012100186005),
    to_complex(- 0.003016982902, - 0.001063857902),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.003001009745, 0.001047884745),
    to_complex(- 0.004159896542, 0.011972396542),
    to_complex(- 0.002985238483, - 0.001032113483),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.002969665021, 0.001016540021),
    to_complex(- 0.004035304858, 0.011847804858),
    to_complex(- 0.002954285372, - 0.001001160372),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.002939095658, 0.000985970658),
    to_complex(- 0.003913783367, 0.011726283367),
    to_complex(- 0.002924092100, - 0.000970967100),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.002909271021, 0.000956146021),
    to_complex(- 0.003795211147, 0.011607711147),
    to_complex(- 0.002894628836, - 0.000941503836),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.002880162056, 0.000927037056),
    to_complex(- 0.003679473509, 0.011491973509),
    to_complex(- 0.002865867281, - 0.000912742281),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.002851741196, 0.000898616196),
    to_complex(- 0.003566461600, 0.011378961600),
    to_complex(- 0.002837780572, - 0.000884655572),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.002823982260, 0.000870857260),
    to_complex(- 0.003456072034, 0.011268572034),
    to_complex(- 0.002810343190, - 0.000857218190),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.002796860370, 0.000843735370),
    to_complex(- 0.003348206556, 0.011160706556),
    to_complex(- 0.002783530881, - 0.000830405881),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.002770351874, 0.000817226874),
    to_complex(- 0.003242771724, 0.011055271724),
    to_complex(- 0.002757320572, - 0.000804195572),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.002744434265, 0.000791309265),
    to_complex(- 0.003139678618, 0.010952178618),
    to_complex(- 0.002731690306, - 0.000778565306),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.002719086115, 0.000765961115),
    to_complex(- 0.003038842571, 0.010851342571),
    to_complex(- 0.002706619172, - 0.000753494172),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.002694287015, 0.000741162015),
    to_complex(- 0.002940182915, 0.010752682915),
    to_complex(- 0.002682087243, - 0.000728962243),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.002670017508, 0.000716892508),
    to_complex(- 0.002843622748, 0.010656122748),
    to_complex(- 0.002658075520, - 0.000704950520),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.002646259040, 0.000693134040),
    to_complex(- 0.002749088717, 0.010561588717),
    to_complex(- 0.002634565879, - 0.000681440879),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.002622993902, 0.000669868902),
    to_complex(- 0.002656510811, 0.010469010811),
    to_complex(- 0.002611541020, - 0.000658416020),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.002600205190, 0.000647080190),
    to_complex(- 0.002565822181, 0.010378322181),
    to_complex(- 0.002588984419, - 0.000635859419),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.002577876754, 0.000624751754),
    to_complex(- 0.002476958953, 0.010289458953),
    to_complex(- 0.002566880288, - 0.000613755288),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.002555993155, 0.000602868155),
    to_complex(- 0.002389860070, 0.010202360070),
    to_complex(- 0.002545213532, - 0.000592088532),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.002534539634, 0.000581414634),
    to_complex(- 0.002304467136, 0.010116967136),
    to_complex(- 0.002523969714, - 0.000570844714),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.002513502065, 0.000560377065),
    to_complex(- 0.002220724273, 0.010033224273),
    to_complex(- 0.002503135015, - 0.000550010015),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.002492866930, 0.000539741930),
    to_complex(- 0.002138577986, 0.009951077986),
    to_complex(- 0.002482696207, - 0.000529571207),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.002472621279, 0.000519496279),
    to_complex(- 0.002057977034, 0.009870477034),
    to_complex(- 0.002462640614, - 0.000509515614),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.002452752708, 0.000499627708),
    to_complex(- 0.001978872317, 0.009791372317),
    to_complex(- 0.002442956091, - 0.000489831091),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.002433249323, 0.000480124323),
    to_complex(- 0.001901216762, 0.009713716762),
    to_complex(- 0.002423630993, - 0.000470505993),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.002414099720, 0.000460974720),
    to_complex(- 0.001824965219, 0.009637465219),
    to_complex(- 0.002404654149, - 0.000451529149),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.002395292954, 0.000442167954),
    to_complex(- 0.001750074363, 0.009562574363),
    to_complex(- 0.002386014836, - 0.000432889836),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.002376818523, 0.000423693523),
    to_complex(- 0.001676502604, 0.009489002604),
    to_complex(- 0.002367702764, - 0.000414577764),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.002358666339, 0.000405541339),
    to_complex(- 0.001604209999, 0.009416709999),
    to_complex(- 0.002349708046, - 0.000396583046),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.002340826712, 0.000387701712),
    to_complex(- 0.001533158172, 0.009345658172),
    to_complex(- 0.002332021183, - 0.000378896183),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.002323290330, 0.000370165330),
    to_complex(- 0.001463310237, 0.009275810237),
    to_complex(- 0.002314633044, - 0.000361508044),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.002306048238, 0.000352923238),
    to_complex(- 0.001394630723, 0.009207130723),
    to_complex(- 0.002297534846, - 0.000344409846),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.002289091823, 0.000335966823),
    to_complex(- 0.001327085514, 0.009139585514),
    to_complex(- 0.002280718143, - 0.000327593143),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.002272412799, 0.000319287799),
    to_complex(- 0.001260641774, 0.009073141774),
    to_complex(- 0.002264174804, - 0.000311049804),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.002256003188, 0.000302878188),
    to_complex(- 0.001195267898, 0.009007767898),
    to_complex(- 0.002247897001, - 0.000294772001),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.002239855309, 0.000286730309),
    to_complex(- 0.001130933446, 0.008943433446),
    to_complex(- 0.002231877196, - 0.000278752196),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.002223961762, 0.000270836762),
    to_complex(- 0.001067609092, 0.008880109092),
    to_complex(- 0.002216108124, - 0.000262983124),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.002208315416, 0.000255190416),
    to_complex(- 0.001005266576, 0.008817766576),
    to_complex(- 0.002200582786, - 0.000247457786),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.002192909398, 0.000239784398),
    to_complex(- 0.000943878651, 0.008756378651),
    to_complex(- 0.002185294431, - 0.000232169431),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.002177737079, 0.000224612079),
    to_complex(- 0.000883419041, 0.008695919041),
    to_complex(- 0.002170236549, - 0.000217111549),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.002162792064, 0.000209667064),
    to_complex(- 0.000823862396, 0.008636362396),
    to_complex(- 0.002155402859, - 0.000202277859),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.002148068183, 0.000194943183),
    to_complex(- 0.000765184251, 0.008577684251),
    to_complex(- 0.002140787299, - 0.000187662299),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.002133559480, 0.000180434480),
    to_complex(- 0.000707360990, 0.008519860990),
    to_complex(- 0.002126384015, - 0.000173259015),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.002119260203, 0.000166135203),
    to_complex(- 0.000650369804, 0.008462869804),
    to_complex(- 0.002112187355, - 0.000159062355),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.002105164796, 0.000152039796),
    to_complex(- 0.000594188662, 0.008406688662),
    to_complex(- 0.002098191859, - 0.000145066859),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.002091267891, 0.000138142891),
    to_complex(- 0.000538796274, 0.008351296274),
    to_complex(- 0.002084392248, - 0.000131267248),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.002077564299, 0.000124439299),
    to_complex(- 0.000484172060, 0.008296672060),
    to_complex(- 0.002070783422, - 0.000117658422),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.002064049005, 0.000110924005),
    to_complex(- 0.000430296122, 0.008242796122),
    to_complex(- 0.002057360447, - 0.000104235447),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.002050717156, 0.000097592156),
    to_complex(- 0.000377149215, 0.008189649215),
    to_complex(- 0.002044118551, - 0.000090993551),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.002037564059, 0.000084439059),
    to_complex(- 0.000324712718, 0.008137212718),
    to_complex(- 0.002031053118, - 0.000077928118),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.002024585173, 0.000071460173),
    to_complex(- 0.000272968613, 0.008085468613),
    to_complex(- 0.002018159679, - 0.000065034679),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.002011776100, 0.000058651100),
    to_complex(- 0.000221899454, 0.008034399454),
    to_complex(- 0.002005433908, - 0.000052308908),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001999132584, 0.000046007584),
    to_complex(- 0.000171488351, 0.007983988351),
    to_complex(- 0.001992871617, - 0.000039746617),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001986650503, 0.000033525503),
    to_complex(- 0.000121718942, 0.007934218942),
    to_complex(- 0.001980468746, - 0.000027343746),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001974325860, 0.000021200860),
    to_complex(- 0.000072575374, 0.007885075374),
    to_complex(- 0.001968221365, - 0.000015096365),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001962154787, 0.000009029787),
    to_complex(- 0.000024042286, 0.007836542286),
    to_complex(- 0.001956125662, - 0.000003000662),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001950133530, - 0.000002991470),
    to_complex(0.000023895215, 0.007788604785),
    to_complex(- 0.001944177942, 0.000008947058),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001938258452, - 0.000014866548),
    to_complex(0.000071251570, 0.007741248430),
    to_complex(- 0.001932374624, 0.000020750376),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001926526025, - 0.000026598975),
    to_complex(0.000118040785, 0.007694459215),
    to_complex(- 0.001920712231, 0.000032412769),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001914932825, - 0.000038192175),
    to_complex(0.000164276448, 0.007648223552),
    to_complex(- 0.001909187394, 0.000043937606),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001903475532, - 0.000049649468),
    to_complex(0.000209971745, 0.007602528255),
    to_complex(- 0.001897796839, 0.000055328161),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001892150921, - 0.000060974079),
    to_complex(0.000255139475, 0.007557360525),
    to_complex(- 0.001886537390, 0.000066587610),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001880955863, - 0.000072169137),
    to_complex(0.000299792066, 0.007512707934),
    to_complex(- 0.001875405964, 0.000077719036),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001869887319, - 0.000083237681),
    to_complex(0.000343941586, 0.007468558414),
    to_complex(- 0.001864399564, 0.000088725436),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001858942337, - 0.000094182663),
    to_complex(0.000387599758, 0.007424900242),
    to_complex(- 0.001853515283, 0.000099609717),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001848118049, - 0.000105006951),
    to_complex(0.000430777971, 0.007381722029),
    to_complex(- 0.001842750291, 0.000110374709),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001837411667, - 0.000115713333),
    to_complex(0.000473487297, 0.007339012703),
    to_complex(- 0.001832101842, 0.000121023158),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001826820483, - 0.000126304517),
    to_complex(0.000515738495, 0.007296761505),
    to_complex(- 0.001821567264, 0.000131557736),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001816341862, - 0.000136783138),
    to_complex(0.000557542028, 0.007254957972),
    to_complex(- 0.001811143959, 0.000141981041),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001805973242, - 0.000147151758),
    to_complex(0.000598908073, 0.007213591927),
    to_complex(- 0.001800829402, 0.000152295598),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001795712133, - 0.000157412867),
    to_complex(0.000639846527, 0.007172653473),
    to_complex(- 0.001790621134, 0.000162503866),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001785556109, - 0.000167568891),
    to_complex(0.000680367022, 0.007132132978),
    to_complex(- 0.001780516764, 0.000172608236),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001775502811, - 0.000177622189),
    to_complex(0.000720478930, 0.007092021070),
    to_complex(- 0.001770513965, 0.000182611035),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001765549944, - 0.000187575056),
    to_complex(0.000760191377, 0.007052308623),
    to_complex(- 0.001760610470, 0.000192514530),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001755695270, - 0.000197429730),
    to_complex(0.000799513246, 0.007012986754),
    to_complex(- 0.001750804074, 0.000202320926),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001745936614, - 0.000207188386),
    to_complex(0.000838453189, 0.006974046811),
    to_complex(- 0.001741092627, 0.000212032373),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001736271854, - 0.000216853146),
    to_complex(0.000877019632, 0.006935480368),
    to_complex(- 0.001731474037, 0.000221650963),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001726698924, - 0.000226426076),
    to_complex(0.000915220787, 0.006897279213),
    to_complex(- 0.001721946264, 0.000231178736),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001717215811, - 0.000235909189),
    to_complex(0.000953064656, 0.006859435344),
    to_complex(- 0.001712507321, 0.000240617679),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001707820553, - 0.000245304447),
    to_complex(0.000990559037, 0.006821940963),
    to_complex(- 0.001703155270, 0.000249969730),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001698511237, - 0.000254613763),
    to_complex(0.001027711535, 0.006784788465),
    to_complex(- 0.001693888222, 0.000259236778),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001689285997, - 0.000263839003),
    to_complex(0.001064529563, 0.006747970437),
    to_complex(- 0.001684704335, 0.000268420665),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001680143014, - 0.000272981986),
    to_complex(0.001101020354, 0.006711479646),
    to_complex(- 0.001675601812, 0.000277523188),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001671080513, - 0.000282044487),
    to_complex(0.001137190962, 0.006675309038),
    to_complex(- 0.001666578901, 0.000286546099),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001662096763, - 0.000291028237),
    to_complex(0.001173048272, 0.006639451728),
    to_complex(- 0.001657633891, 0.000295491109),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001653190075, - 0.000299934925),
    to_complex(0.001208599002, 0.006603900998),
    to_complex(- 0.001648765112, 0.000304359888),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001644358798, - 0.000308766202),
    to_complex(0.001243849710, 0.006568650290),
    to_complex(- 0.001639970935, 0.000313154065),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001635601323, - 0.000317523677),
    to_complex(0.001278806799, 0.006533693201),
    to_complex(- 0.001631249768, 0.000321875232),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001626916076, - 0.000326208924),
    to_complex(0.001313476521, 0.006499023479),
    to_complex(- 0.001622600057, 0.000330524943),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001618301523, - 0.000334823477),
    to_complex(0.001347864986, 0.006464635014),
    to_complex(- 0.001614020285, 0.000339104715),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001609756162, - 0.000343368838),
    to_complex(0.001381978160, 0.006430521840),
    to_complex(- 0.001605508969, 0.000347616031),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001601278527, - 0.000351846473),
    to_complex(0.001415821873, 0.006396678127),
    to_complex(- 0.001597064658, 0.000356060342),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001592867186, - 0.000360257814),
    to_complex(0.001449401825, 0.006363098175),
    to_complex(- 0.001588685936, 0.000364439064),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001584520737, - 0.000368604263),
    to_complex(0.001482723586, 0.006329776414),
    to_complex(- 0.001580371419, 0.000372753581),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001576237813, - 0.000376887187),
    to_complex(0.001515792602, 0.006296707398),
    to_complex(- 0.001572119752, 0.000381005248),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001568017072, - 0.000385107928),
    to_complex(0.001548614202, 0.006263885798),
    to_complex(- 0.001563929611, 0.000389195389),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001559857207, - 0.000393267793),
    to_complex(0.001581193595, 0.006231306405),
    to_complex(- 0.001555799701, 0.000397325299),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001551756935, - 0.000401368065),
    to_complex(0.001613535878, 0.006198964122),
    to_complex(- 0.001547728753, 0.000405396247),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001543715002, - 0.000409409998),
    to_complex(0.001645646040, 0.006166853960),
    to_complex(- 0.001539715528, 0.000413409472),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001535730182, - 0.000417394818),
    to_complex(0.001677528964, 0.006134971036),
    to_complex(- 0.001531758812, 0.000421366188),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001527801273, - 0.000425323727),
    to_complex(0.001709189427, 0.006103310573),
    to_complex(- 0.001523857416, 0.000429267584),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001519927099, - 0.000433197901),
    to_complex(0.001740632111, 0.006071867889),
    to_complex(- 0.001516010177, 0.000437114823),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001512106509, - 0.000441018491),
    to_complex(0.001771861597, 0.006040638403),
    to_complex(- 0.001508215954, 0.000444909046),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001504338374, - 0.000448786626),
    to_complex(0.001802882374, 0.006009617626),
    to_complex(- 0.001500473631, 0.000452651369),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001496621590, - 0.000456503410),
    to_complex(0.001833698841, 0.005978801159),
    to_complex(- 0.001492782115, 0.000460342885),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001488955073, - 0.000464169927),
    to_complex(0.001864315308, 0.005948184692),
    to_complex(- 0.001485140332, 0.000467984668),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001481337762, - 0.000471787238),
    to_complex(0.001894735997, 0.005917764003),
    to_complex(- 0.001477547233, 0.000475577767),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001473768618, - 0.000479356382),
    to_complex(0.001924965050, 0.005887534950),
    to_complex(- 0.001470001788, 0.000483123212),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001466246619, - 0.000486878381),
    to_complex(0.001955006527, 0.005857493473),
    to_complex(- 0.001462502986, 0.000490622014),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001458770766, - 0.000494354234),
    to_complex(0.001984864410, 0.005827635590),
    to_complex(- 0.001455049837, 0.000498075163),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001451340077, - 0.000501784923),
    to_complex(0.002014542605, 0.005797957395),
    to_complex(- 0.001447641368, 0.000505483632),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001443953590, - 0.000509171410),
    to_complex(0.002044044943, 0.005768455057),
    to_complex(- 0.001440276627, 0.000512848373),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001436610361, - 0.000516514639),
    to_complex(0.002073375186, 0.005739124814),
    to_complex(- 0.001432954677, 0.000520170323),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001429309462, - 0.000523815538),
    to_complex(0.002102537023, 0.005709962977),
    to_complex(- 0.001425674601, 0.000527450399),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001422049983, - 0.000531075017),
    to_complex(0.002131534078, 0.005680965922),
    to_complex(- 0.001418435497, 0.000534689503),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001414831031, - 0.000538293969),
    to_complex(0.002160369910, 0.005652130090),
    to_complex(- 0.001411236478, 0.000541888522),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001407651729, - 0.000545473271),
    to_complex(0.002189048012, 0.005623451988),
    to_complex(- 0.001404076676, 0.000549048324),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001400511213, - 0.000552613787),
    to_complex(0.002217571818, 0.005594928182),
    to_complex(- 0.001396955236, 0.000556169764),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001393408639, - 0.000559716361),
    to_complex(0.002245944699, 0.005566555301),
    to_complex(- 0.001389871318, 0.000563253682),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001386343172, - 0.000566781828),
    to_complex(0.002274169970, 0.005538330030),
    to_complex(- 0.001382824098, 0.000570300902),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001379313996, - 0.000573811004),
    to_complex(0.002302250889, 0.005510249111),
    to_complex(- 0.001375812765, 0.000577312235),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001372320306, - 0.000580804694),
    to_complex(0.002330190659, 0.005482309341),
    to_complex(- 0.001368836521, 0.000584288479),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001365361311, - 0.000587763689),
    to_complex(0.002357992430, 0.005454507570),
    to_complex(- 0.001361894581, 0.000591230419),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001358436235, - 0.000594688765),
    to_complex(0.002385659299, 0.005426840701),
    to_complex(- 0.001354986176, 0.000598138824),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001351544311, - 0.000601580689),
    to_complex(0.002413194315, 0.005399305685),
    to_complex(- 0.001348110545, 0.000605014455),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001344684786, - 0.000608440214),
    to_complex(0.002440600477, 0.005371899523),
    to_complex(- 0.001341266942, 0.000611858058),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001337856921, - 0.000615268079),
    to_complex(0.002467880736, 0.005344619264),
    to_complex(- 0.001334454633, 0.000618670367),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001331059986, - 0.000622065014),
    to_complex(0.002495037998, 0.005317462002),
    to_complex(- 0.001327672892, 0.000625452108),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001324293262, - 0.000628831738),
    to_complex(0.002522075124, 0.005290424876),
    to_complex(- 0.001320921008, 0.000632203992),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001317556043, - 0.000635568957),
    to_complex(0.002548994933, 0.005263505067),
    to_complex(- 0.001314198280, 0.000638926720),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001310847632, - 0.000642277368),
    to_complex(0.002575800200, 0.005236699800),
    to_complex(- 0.001307504015, 0.000645620985),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001304167343, - 0.000648957657),
    to_complex(0.002602493661, 0.005210006339),
    to_complex(- 0.001300837532, 0.000652287468),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001297514499, - 0.000655610501),
    to_complex(0.002629078010, 0.005183421990),
    to_complex(- 0.001294198160, 0.000658926840),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001290888433, - 0.000662236567),
    to_complex(0.002655555906, 0.005156944094),
    to_complex(- 0.001287585236, 0.000665539764),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001284288489, - 0.000668836511),
    to_complex(0.002681929968, 0.005130570032),
    to_complex(- 0.001280998109, 0.000672126891),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001277714017, - 0.000675410983),
    to_complex(0.002708202781, 0.005104297219),
    to_complex(- 0.001274436134, 0.000678688866),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001271164380, - 0.000681960620),
    to_complex(0.002734376894, 0.005078123106),
    to_complex(- 0.001267898676, 0.000685226324),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001264638945, - 0.000688486055),
    to_complex(0.002760454821, 0.005052045179),
    to_complex(- 0.001261385109, 0.000691739891),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001258137090, - 0.000694987910),
    to_complex(0.002786439045, 0.005026060955),
    to_complex(- 0.001254894813, 0.000698230187),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001251658201, - 0.000701466799),
    to_complex(0.002812332016, 0.005000167984),
    to_complex(- 0.001248427179, 0.000704697821),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001245201671, - 0.000707923329),
    to_complex(0.002838136153, 0.004974363847),
    to_complex(- 0.001241981603, 0.000711143397),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001238766901, - 0.000714358099),
    to_complex(0.002863853847, 0.004948646153),
    to_complex(- 0.001235557490, 0.000717567510),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001232353298, - 0.000720771702),
    to_complex(0.002889487457, 0.004923012543),
    to_complex(- 0.001229154251, 0.000723970749),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001225960278, - 0.000727164722),
    to_complex(0.002915039317, 0.004897460683),
    to_complex(- 0.001222771305, 0.000730353695),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001219587262, - 0.000733537738),
    to_complex(0.002940511731, 0.004871988269),
    to_complex(- 0.001216408078, 0.000736716922),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001213233680, - 0.000739891320),
    to_complex(0.002965906980, 0.004846593020),
    to_complex(- 0.001210064000, 0.000743061000),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001206898967, - 0.000746226033),
    to_complex(0.002991227316, 0.004821272684),
    to_complex(- 0.001203738511, 0.000749386489),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001200582563, - 0.000752542437),
    to_complex(0.003016474969, 0.004796025031),
    to_complex(- 0.001197431054, 0.000755693946),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001194283916, - 0.000758841084),
    to_complex(0.003041652144, 0.004770847856),
    to_complex(- 0.001191141079, 0.000761983921),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001188002478, - 0.000765122522),
    to_complex(0.003066761025, 0.004745738975),
    to_complex(- 0.001184868043, 0.000768256957),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001181737708, - 0.000771387292),
    to_complex(0.003091803772, 0.004720696228),
    to_complex(- 0.001178611406, 0.000774513594),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001175489070, - 0.000777635930),
    to_complex(0.003116782524, 0.004695717476),
    to_complex(- 0.001172370635, 0.000780754365),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001169256033, - 0.000783868967),
    to_complex(0.003141699400, 0.004670800600),
    to_complex(- 0.001166145201, 0.000786979799),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001163038071, - 0.000790086929),
    to_complex(0.003166556499, 0.004645943501),
    to_complex(- 0.001159934581, 0.000793190419),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001156834663, - 0.000796290337),
    to_complex(0.003191355901, 0.004621144099),
    to_complex(- 0.001153738255, 0.000799386745),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001150645292, - 0.000802479708),
    to_complex(0.003216099668, 0.004596400332),
    to_complex(- 0.001147555711, 0.000805569289),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001144469447, - 0.000808655553),
    to_complex(0.003240789843, 0.004571710157),
    to_complex(- 0.001141386437, 0.000811738563),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001138306619, - 0.000814818381),
    to_complex(0.003265428455, 0.004547071545),
    to_complex(- 0.001135229928, 0.000817895072),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001132156304, - 0.000820968696),
    to_complex(0.003290017513, 0.004522482487),
    to_complex(- 0.001129085683, 0.000824039317),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001126018003, - 0.000827106997),
    to_complex(0.003314559013, 0.004497940987),
    to_complex(- 0.001122953203, 0.000830171797),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001119891220, - 0.000833233780),
    to_complex(0.003339054936, 0.004473445064),
    to_complex(- 0.001116831993, 0.000836293007),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001113775462, - 0.000839349538),
    to_complex(0.003363507249, 0.004448992751),
    to_complex(- 0.001110721565, 0.000842403435),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001107670240, - 0.000845454760),
    to_complex(0.003387917903, 0.004424582097),
    to_complex(- 0.001104621429, 0.000848503571),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001101575069, - 0.000851549931),
    to_complex(0.003412288839, 0.004400211161),
    to_complex(- 0.001098531102, 0.000854593898),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001095489466, - 0.000857635534),
    to_complex(0.003436621984, 0.004375878016),
    to_complex(- 0.001092450102, 0.000860674898),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001089412951, - 0.000863712049),
    to_complex(0.003460919255, 0.004351580745),
    to_complex(- 0.001086377952, 0.000866747048),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001083345047, - 0.000869779953),
    to_complex(0.003485182556, 0.004327317444),
    to_complex(- 0.001080314176, 0.000872810824),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001077285280, - 0.000875839720),
    to_complex(0.003509413782, 0.004303086218),
    to_complex(- 0.001074258301, 0.000878866699),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001071233179, - 0.000881891821),
    to_complex(0.003533614817, 0.004278885183),
    to_complex(- 0.001068209855, 0.000884915145),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001065188273, - 0.000887936727),
    to_complex(0.003557787537, 0.004254712463),
    to_complex(- 0.001062168372, 0.000890956628),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001059150095, - 0.000893974905),
    to_complex(0.003581933809, 0.004230566191),
    to_complex(- 0.001056133384, 0.000896991616),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001053118181, - 0.000900006819),
    to_complex(0.003606055491, 0.004206444509),
    to_complex(- 0.001050104428, 0.000903020572),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001047092068, - 0.000906032932),
    to_complex(0.003630154434, 0.004182345566),
    to_complex(- 0.001044081042, 0.000909043958),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001041071293, - 0.000912053707),
    to_complex(0.003654232484, 0.004158267516),
    to_complex(- 0.001038062763, 0.000915062237),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001035055396, - 0.000918069604),
    to_complex(0.003678291477, 0.004134208523),
    to_complex(- 0.001032049134, 0.000921075866),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001029043920, - 0.000924081080),
    to_complex(0.003702333246, 0.004110166754),
    to_complex(- 0.001026039697, 0.000927085303),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001023036408, - 0.000930088592),
    to_complex(0.003726359619, 0.004086140381),
    to_complex(- 0.001020033995, 0.000933091005),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001017032402, - 0.000936092598),
    to_complex(0.003750372416, 0.004062127584),
    to_complex(- 0.001014031573, 0.000939093427),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001011031450, - 0.000942093550),
    to_complex(0.003774373458, 0.004038126542),
    to_complex(- 0.001008031977, 0.000945093023),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.001005033096, - 0.000948091904),
    to_complex(0.003798364557, 0.004014135443),
    to_complex(- 0.001002034752, 0.000951090248),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000999036888, - 0.000954088112),
    to_complex(0.003822347526, 0.003990152474),
    to_complex(- 0.000996039447, 0.000957085553),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000993042373, - 0.000960082627),
    to_complex(0.003846324175, 0.003966175825),
    to_complex(- 0.000990045610, 0.000963079390),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000987049100, - 0.000966075900),
    to_complex(0.003870296310, 0.003942203690),
    to_complex(- 0.000984052787, 0.000969072213),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000981056616, - 0.000972068384),
    to_complex(0.003894265737, 0.003918234263),
    to_complex(- 0.000978060529, 0.000975064471),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000975064471, - 0.000978060529),
    to_complex(0.003918234263, 0.003894265737),
    to_complex(- 0.000972068384, 0.000981056616),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000969072213, - 0.000984052787),
    to_complex(0.003942203690, 0.003870296310),
    to_complex(- 0.000966075900, 0.000987049100),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000963079390, - 0.000990045610),
    to_complex(0.003966175825, 0.003846324175),
    to_complex(- 0.000960082627, 0.000993042373),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000957085553, - 0.000996039447),
    to_complex(0.003990152474, 0.003822347526),
    to_complex(- 0.000954088112, 0.000999036888),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000951090248, - 0.001002034752),
    to_complex(0.004014135443, 0.003798364557),
    to_complex(- 0.000948091904, 0.001005033096),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000945093023, - 0.001008031977),
    to_complex(0.004038126542, 0.003774373458),
    to_complex(- 0.000942093550, 0.001011031450),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000939093427, - 0.001014031573),
    to_complex(0.004062127584, 0.003750372416),
    to_complex(- 0.000936092598, 0.001017032402),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000933091005, - 0.001020033995),
    to_complex(0.004086140381, 0.003726359619),
    to_complex(- 0.000930088592, 0.001023036408),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000927085303, - 0.001026039697),
    to_complex(0.004110166754, 0.003702333246),
    to_complex(- 0.000924081080, 0.001029043920),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000921075866, - 0.001032049134),
    to_complex(0.004134208523, 0.003678291477),
    to_complex(- 0.000918069604, 0.001035055396),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000915062237, - 0.001038062763),
    to_complex(0.004158267516, 0.003654232484),
    to_complex(- 0.000912053707, 0.001041071293),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000909043958, - 0.001044081042),
    to_complex(0.004182345566, 0.003630154434),
    to_complex(- 0.000906032932, 0.001047092068),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000903020572, - 0.001050104428),
    to_complex(0.004206444509, 0.003606055491),
    to_complex(- 0.000900006819, 0.001053118181),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000896991616, - 0.001056133384),
    to_complex(0.004230566191, 0.003581933809),
    to_complex(- 0.000893974905, 0.001059150095),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000890956628, - 0.001062168372),
    to_complex(0.004254712463, 0.003557787537),
    to_complex(- 0.000887936727, 0.001065188273),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000884915145, - 0.001068209855),
    to_complex(0.004278885183, 0.003533614817),
    to_complex(- 0.000881891821, 0.001071233179),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000878866699, - 0.001074258301),
    to_complex(0.004303086218, 0.003509413782),
    to_complex(- 0.000875839720, 0.001077285280),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000872810824, - 0.001080314176),
    to_complex(0.004327317444, 0.003485182556),
    to_complex(- 0.000869779953, 0.001083345047),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000866747048, - 0.001086377952),
    to_complex(0.004351580745, 0.003460919255),
    to_complex(- 0.000863712049, 0.001089412951),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000860674898, - 0.001092450102),
    to_complex(0.004375878016, 0.003436621984),
    to_complex(- 0.000857635534, 0.001095489466),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000854593898, - 0.001098531102),
    to_complex(0.004400211161, 0.003412288839),
    to_complex(- 0.000851549931, 0.001101575069),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000848503571, - 0.001104621429),
    to_complex(0.004424582097, 0.003387917903),
    to_complex(- 0.000845454760, 0.001107670240),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000842403435, - 0.001110721565),
    to_complex(0.004448992751, 0.003363507249),
    to_complex(- 0.000839349538, 0.001113775462),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000836293007, - 0.001116831993),
    to_complex(0.004473445064, 0.003339054936),
    to_complex(- 0.000833233780, 0.001119891220),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000830171797, - 0.001122953203),
    to_complex(0.004497940987, 0.003314559013),
    to_complex(- 0.000827106997, 0.001126018003),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000824039317, - 0.001129085683),
    to_complex(0.004522482487, 0.003290017513),
    to_complex(- 0.000820968696, 0.001132156304),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000817895072, - 0.001135229928),
    to_complex(0.004547071545, 0.003265428455),
    to_complex(- 0.000814818381, 0.001138306619),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000811738563, - 0.001141386437),
    to_complex(0.004571710157, 0.003240789843),
    to_complex(- 0.000808655553, 0.001144469447),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000805569289, - 0.001147555711),
    to_complex(0.004596400332, 0.003216099668),
    to_complex(- 0.000802479708, 0.001150645292),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000799386745, - 0.001153738255),
    to_complex(0.004621144099, 0.003191355901),
    to_complex(- 0.000796290337, 0.001156834663),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000793190419, - 0.001159934581),
    to_complex(0.004645943501, 0.003166556499),
    to_complex(- 0.000790086929, 0.001163038071),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000786979799, - 0.001166145201),
    to_complex(0.004670800600, 0.003141699400),
    to_complex(- 0.000783868967, 0.001169256033),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000780754365, - 0.001172370635),
    to_complex(0.004695717476, 0.003116782524),
    to_complex(- 0.000777635930, 0.001175489070),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000774513594, - 0.001178611406),
    to_complex(0.004720696228, 0.003091803772),
    to_complex(- 0.000771387292, 0.001181737708),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000768256957, - 0.001184868043),
    to_complex(0.004745738975, 0.003066761025),
    to_complex(- 0.000765122522, 0.001188002478),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000761983921, - 0.001191141079),
    to_complex(0.004770847856, 0.003041652144),
    to_complex(- 0.000758841084, 0.001194283916),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000755693946, - 0.001197431054),
    to_complex(0.004796025031, 0.003016474969),
    to_complex(- 0.000752542437, 0.001200582563),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000749386489, - 0.001203738511),
    to_complex(0.004821272684, 0.002991227316),
    to_complex(- 0.000746226033, 0.001206898967),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000743061000, - 0.001210064000),
    to_complex(0.004846593020, 0.002965906980),
    to_complex(- 0.000739891320, 0.001213233680),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000736716922, - 0.001216408078),
    to_complex(0.004871988269, 0.002940511731),
    to_complex(- 0.000733537738, 0.001219587262),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000730353695, - 0.001222771305),
    to_complex(0.004897460683, 0.002915039317),
    to_complex(- 0.000727164722, 0.001225960278),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000723970749, - 0.001229154251),
    to_complex(0.004923012543, 0.002889487457),
    to_complex(- 0.000720771702, 0.001232353298),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000717567510, - 0.001235557490),
    to_complex(0.004948646153, 0.002863853847),
    to_complex(- 0.000714358099, 0.001238766901),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000711143397, - 0.001241981603),
    to_complex(0.004974363847, 0.002838136153),
    to_complex(- 0.000707923329, 0.001245201671),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000704697821, - 0.001248427179),
    to_complex(0.005000167984, 0.002812332016),
    to_complex(- 0.000701466799, 0.001251658201),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000698230187, - 0.001254894813),
    to_complex(0.005026060955, 0.002786439045),
    to_complex(- 0.000694987910, 0.001258137090),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000691739891, - 0.001261385109),
    to_complex(0.005052045179, 0.002760454821),
    to_complex(- 0.000688486055, 0.001264638945),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000685226324, - 0.001267898676),
    to_complex(0.005078123106, 0.002734376894),
    to_complex(- 0.000681960620, 0.001271164380),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000678688866, - 0.001274436134),
    to_complex(0.005104297219, 0.002708202781),
    to_complex(- 0.000675410983, 0.001277714017),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000672126891, - 0.001280998109),
    to_complex(0.005130570032, 0.002681929968),
    to_complex(- 0.000668836511, 0.001284288489),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000665539764, - 0.001287585236),
    to_complex(0.005156944094, 0.002655555906),
    to_complex(- 0.000662236567, 0.001290888433),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000658926840, - 0.001294198160),
    to_complex(0.005183421990, 0.002629078010),
    to_complex(- 0.000655610501, 0.001297514499),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000652287468, - 0.001300837532),
    to_complex(0.005210006339, 0.002602493661),
    to_complex(- 0.000648957657, 0.001304167343),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000645620985, - 0.001307504015),
    to_complex(0.005236699800, 0.002575800200),
    to_complex(- 0.000642277368, 0.001310847632),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000638926720, - 0.001314198280),
    to_complex(0.005263505067, 0.002548994933),
    to_complex(- 0.000635568957, 0.001317556043),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000632203992, - 0.001320921008),
    to_complex(0.005290424876, 0.002522075124),
    to_complex(- 0.000628831738, 0.001324293262),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000625452108, - 0.001327672892),
    to_complex(0.005317462002, 0.002495037998),
    to_complex(- 0.000622065014, 0.001331059986),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000618670367, - 0.001334454633),
    to_complex(0.005344619264, 0.002467880736),
    to_complex(- 0.000615268079, 0.001337856921),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000611858058, - 0.001341266942),
    to_complex(0.005371899523, 0.002440600477),
    to_complex(- 0.000608440214, 0.001344684786),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000605014455, - 0.001348110545),
    to_complex(0.005399305685, 0.002413194315),
    to_complex(- 0.000601580689, 0.001351544311),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000598138824, - 0.001354986176),
    to_complex(0.005426840701, 0.002385659299),
    to_complex(- 0.000594688765, 0.001358436235),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000591230419, - 0.001361894581),
    to_complex(0.005454507570, 0.002357992430),
    to_complex(- 0.000587763689, 0.001365361311),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000584288479, - 0.001368836521),
    to_complex(0.005482309341, 0.002330190659),
    to_complex(- 0.000580804694, 0.001372320306),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000577312235, - 0.001375812765),
    to_complex(0.005510249111, 0.002302250889),
    to_complex(- 0.000573811004, 0.001379313996),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000570300902, - 0.001382824098),
    to_complex(0.005538330030, 0.002274169970),
    to_complex(- 0.000566781828, 0.001386343172),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000563253682, - 0.001389871318),
    to_complex(0.005566555301, 0.002245944699),
    to_complex(- 0.000559716361, 0.001393408639),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000556169764, - 0.001396955236),
    to_complex(0.005594928182, 0.002217571818),
    to_complex(- 0.000552613787, 0.001400511213),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000549048324, - 0.001404076676),
    to_complex(0.005623451988, 0.002189048012),
    to_complex(- 0.000545473271, 0.001407651729),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000541888522, - 0.001411236478),
    to_complex(0.005652130090, 0.002160369910),
    to_complex(- 0.000538293969, 0.001414831031),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000534689503, - 0.001418435497),
    to_complex(0.005680965922, 0.002131534078),
    to_complex(- 0.000531075017, 0.001422049983),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000527450399, - 0.001425674601),
    to_complex(0.005709962977, 0.002102537023),
    to_complex(- 0.000523815538, 0.001429309462),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000520170323, - 0.001432954677),
    to_complex(0.005739124814, 0.002073375186),
    to_complex(- 0.000516514639, 0.001436610361),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000512848373, - 0.001440276627),
    to_complex(0.005768455057, 0.002044044943),
    to_complex(- 0.000509171410, 0.001443953590),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000505483632, - 0.001447641368),
    to_complex(0.005797957395, 0.002014542605),
    to_complex(- 0.000501784923, 0.001451340077),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000498075163, - 0.001455049837),
    to_complex(0.005827635590, 0.001984864410),
    to_complex(- 0.000494354234, 0.001458770766),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000490622014, - 0.001462502986),
    to_complex(0.005857493473, 0.001955006527),
    to_complex(- 0.000486878381, 0.001466246619),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000483123212, - 0.001470001788),
    to_complex(0.005887534950, 0.001924965050),
    to_complex(- 0.000479356382, 0.001473768618),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000475577767, - 0.001477547233),
    to_complex(0.005917764003, 0.001894735997),
    to_complex(- 0.000471787238, 0.001481337762),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000467984668, - 0.001485140332),
    to_complex(0.005948184692, 0.001864315308),
    to_complex(- 0.000464169927, 0.001488955073),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000460342885, - 0.001492782115),
    to_complex(0.005978801159, 0.001833698841),
    to_complex(- 0.000456503410, 0.001496621590),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000452651369, - 0.001500473631),
    to_complex(0.006009617626, 0.001802882374),
    to_complex(- 0.000448786626, 0.001504338374),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000444909046, - 0.001508215954),
    to_complex(0.006040638403, 0.001771861597),
    to_complex(- 0.000441018491, 0.001512106509),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000437114823, - 0.001516010177),
    to_complex(0.006071867889, 0.001740632111),
    to_complex(- 0.000433197901, 0.001519927099),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000429267584, - 0.001523857416),
    to_complex(0.006103310573, 0.001709189427),
    to_complex(- 0.000425323727, 0.001527801273),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000421366188, - 0.001531758812),
    to_complex(0.006134971036, 0.001677528964),
    to_complex(- 0.000417394818, 0.001535730182),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000413409472, - 0.001539715528),
    to_complex(0.006166853960, 0.001645646040),
    to_complex(- 0.000409409998, 0.001543715002),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000405396247, - 0.001547728753),
    to_complex(0.006198964122, 0.001613535878),
    to_complex(- 0.000401368065, 0.001551756935),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000397325299, - 0.001555799701),
    to_complex(0.006231306405, 0.001581193595),
    to_complex(- 0.000393267793, 0.001559857207),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000389195389, - 0.001563929611),
    to_complex(0.006263885798, 0.001548614202),
    to_complex(- 0.000385107928, 0.001568017072),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000381005248, - 0.001572119752),
    to_complex(0.006296707398, 0.001515792602),
    to_complex(- 0.000376887187, 0.001576237813),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000372753581, - 0.001580371419),
    to_complex(0.006329776414, 0.001482723586),
    to_complex(- 0.000368604263, 0.001584520737),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000364439064, - 0.001588685936),
    to_complex(0.006363098175, 0.001449401825),
    to_complex(- 0.000360257814, 0.001592867186),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000356060342, - 0.001597064658),
    to_complex(0.006396678127, 0.001415821873),
    to_complex(- 0.000351846473, 0.001601278527),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000347616031, - 0.001605508969),
    to_complex(0.006430521840, 0.001381978160),
    to_complex(- 0.000343368838, 0.001609756162),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000339104715, - 0.001614020285),
    to_complex(0.006464635014, 0.001347864986),
    to_complex(- 0.000334823477, 0.001618301523),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000330524943, - 0.001622600057),
    to_complex(0.006499023479, 0.001313476521),
    to_complex(- 0.000326208924, 0.001626916076),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000321875232, - 0.001631249768),
    to_complex(0.006533693201, 0.001278806799),
    to_complex(- 0.000317523677, 0.001635601323),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000313154065, - 0.001639970935),
    to_complex(0.006568650290, 0.001243849710),
    to_complex(- 0.000308766202, 0.001644358798),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000304359888, - 0.001648765112),
    to_complex(0.006603900998, 0.001208599002),
    to_complex(- 0.000299934925, 0.001653190075),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000295491109, - 0.001657633891),
    to_complex(0.006639451728, 0.001173048272),
    to_complex(- 0.000291028237, 0.001662096763),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000286546099, - 0.001666578901),
    to_complex(0.006675309038, 0.001137190962),
    to_complex(- 0.000282044487, 0.001671080513),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000277523188, - 0.001675601812),
    to_complex(0.006711479646, 0.001101020354),
    to_complex(- 0.000272981986, 0.001680143014),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000268420665, - 0.001684704335),
    to_complex(0.006747970437, 0.001064529563),
    to_complex(- 0.000263839003, 0.001689285997),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000259236778, - 0.001693888222),
    to_complex(0.006784788465, 0.001027711535),
    to_complex(- 0.000254613763, 0.001698511237),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000249969730, - 0.001703155270),
    to_complex(0.006821940963, 0.000990559037),
    to_complex(- 0.000245304447, 0.001707820553),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000240617679, - 0.001712507321),
    to_complex(0.006859435344, 0.000953064656),
    to_complex(- 0.000235909189, 0.001717215811),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000231178736, - 0.001721946264),
    to_complex(0.006897279213, 0.000915220787),
    to_complex(- 0.000226426076, 0.001726698924),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000221650963, - 0.001731474037),
    to_complex(0.006935480368, 0.000877019632),
    to_complex(- 0.000216853146, 0.001736271854),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000212032373, - 0.001741092627),
    to_complex(0.006974046811, 0.000838453189),
    to_complex(- 0.000207188386, 0.001745936614),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000202320926, - 0.001750804074),
    to_complex(0.007012986754, 0.000799513246),
    to_complex(- 0.000197429730, 0.001755695270),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000192514530, - 0.001760610470),
    to_complex(0.007052308623, 0.000760191377),
    to_complex(- 0.000187575056, 0.001765549944),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000182611035, - 0.001770513965),
    to_complex(0.007092021070, 0.000720478930),
    to_complex(- 0.000177622189, 0.001775502811),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000172608236, - 0.001780516764),
    to_complex(0.007132132978, 0.000680367022),
    to_complex(- 0.000167568891, 0.001785556109),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000162503866, - 0.001790621134),
    to_complex(0.007172653473, 0.000639846527),
    to_complex(- 0.000157412867, 0.001795712133),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000152295598, - 0.001800829402),
    to_complex(0.007213591927, 0.000598908073),
    to_complex(- 0.000147151758, 0.001805973242),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000141981041, - 0.001811143959),
    to_complex(0.007254957972, 0.000557542028),
    to_complex(- 0.000136783138, 0.001816341862),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000131557736, - 0.001821567264),
    to_complex(0.007296761505, 0.000515738495),
    to_complex(- 0.000126304517, 0.001826820483),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000121023158, - 0.001832101842),
    to_complex(0.007339012703, 0.000473487297),
    to_complex(- 0.000115713333, 0.001837411667),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000110374709, - 0.001842750291),
    to_complex(0.007381722029, 0.000430777971),
    to_complex(- 0.000105006951, 0.001848118049),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000099609717, - 0.001853515283),
    to_complex(0.007424900242, 0.000387599758),
    to_complex(- 0.000094182663, 0.001858942337),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000088725436, - 0.001864399564),
    to_complex(0.007468558414, 0.000343941586),
    to_complex(- 0.000083237681, 0.001869887319),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000077719036, - 0.001875405964),
    to_complex(0.007512707934, 0.000299792066),
    to_complex(- 0.000072169137, 0.001880955863),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000066587610, - 0.001886537390),
    to_complex(0.007557360525, 0.000255139475),
    to_complex(- 0.000060974079, 0.001892150921),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000055328161, - 0.001897796839),
    to_complex(0.007602528255, 0.000209971745),
    to_complex(- 0.000049649468, 0.001903475532),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000043937606, - 0.001909187394),
    to_complex(0.007648223552, 0.000164276448),
    to_complex(- 0.000038192175, 0.001914932825),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000032412769, - 0.001920712231),
    to_complex(0.007694459215, 0.000118040785),
    to_complex(- 0.000026598975, 0.001926526025),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000020750376, - 0.001932374624),
    to_complex(0.007741248430, 0.000071251570),
    to_complex(- 0.000014866548, 0.001938258452),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.000008947058, - 0.001944177942),
    to_complex(0.007788604785, 0.000023895215),
    to_complex(- 0.000002991470, 0.001950133530),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.000003000662, - 0.001956125662),
    to_complex(0.007836542286, - 0.000024042286),
    to_complex(0.000009029787, 0.001962154787),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.000015096365, - 0.001968221365),
    to_complex(0.007885075374, - 0.000072575374),
    to_complex(0.000021200860, 0.001974325860),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.000027343746, - 0.001980468746),
    to_complex(0.007934218942, - 0.000121718942),
    to_complex(0.000033525503, 0.001986650503),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.000039746617, - 0.001992871617),
    to_complex(0.007983988351, - 0.000171488351),
    to_complex(0.000046007584, 0.001999132584),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.000052308908, - 0.002005433908),
    to_complex(0.008034399454, - 0.000221899454),
    to_complex(0.000058651100, 0.002011776100),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.000065034679, - 0.002018159679),
    to_complex(0.008085468613, - 0.000272968613),
    to_complex(0.000071460173, 0.002024585173),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.000077928118, - 0.002031053118),
    to_complex(0.008137212718, - 0.000324712718),
    to_complex(0.000084439059, 0.002037564059),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.000090993551, - 0.002044118551),
    to_complex(0.008189649215, - 0.000377149215),
    to_complex(0.000097592156, 0.002050717156),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.000104235447, - 0.002057360447),
    to_complex(0.008242796122, - 0.000430296122),
    to_complex(0.000110924005, 0.002064049005),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.000117658422, - 0.002070783422),
    to_complex(0.008296672060, - 0.000484172060),
    to_complex(0.000124439299, 0.002077564299),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.000131267248, - 0.002084392248),
    to_complex(0.008351296274, - 0.000538796274),
    to_complex(0.000138142891, 0.002091267891),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.000145066859, - 0.002098191859),
    to_complex(0.008406688662, - 0.000594188662),
    to_complex(0.000152039796, 0.002105164796),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.000159062355, - 0.002112187355),
    to_complex(0.008462869804, - 0.000650369804),
    to_complex(0.000166135203, 0.002119260203),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.000173259015, - 0.002126384015),
    to_complex(0.008519860990, - 0.000707360990),
    to_complex(0.000180434480, 0.002133559480),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.000187662299, - 0.002140787299),
    to_complex(0.008577684251, - 0.000765184251),
    to_complex(0.000194943183, 0.002148068183),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.000202277859, - 0.002155402859),
    to_complex(0.008636362396, - 0.000823862396),
    to_complex(0.000209667064, 0.002162792064),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.000217111549, - 0.002170236549),
    to_complex(0.008695919041, - 0.000883419041),
    to_complex(0.000224612079, 0.002177737079),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.000232169431, - 0.002185294431),
    to_complex(0.008756378651, - 0.000943878651),
    to_complex(0.000239784398, 0.002192909398),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.000247457786, - 0.002200582786),
    to_complex(0.008817766576, - 0.001005266576),
    to_complex(0.000255190416, 0.002208315416),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.000262983124, - 0.002216108124),
    to_complex(0.008880109092, - 0.001067609092),
    to_complex(0.000270836762, 0.002223961762),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.000278752196, - 0.002231877196),
    to_complex(0.008943433446, - 0.001130933446),
    to_complex(0.000286730309, 0.002239855309),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.000294772001, - 0.002247897001),
    to_complex(0.009007767898, - 0.001195267898),
    to_complex(0.000302878188, 0.002256003188),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.000311049804, - 0.002264174804),
    to_complex(0.009073141774, - 0.001260641774),
    to_complex(0.000319287799, 0.002272412799),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.000327593143, - 0.002280718143),
    to_complex(0.009139585514, - 0.001327085514),
    to_complex(0.000335966823, 0.002289091823),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.000344409846, - 0.002297534846),
    to_complex(0.009207130723, - 0.001394630723),
    to_complex(0.000352923238, 0.002306048238),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.000361508044, - 0.002314633044),
    to_complex(0.009275810237, - 0.001463310237),
    to_complex(0.000370165330, 0.002323290330),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.000378896183, - 0.002332021183),
    to_complex(0.009345658172, - 0.001533158172),
    to_complex(0.000387701712, 0.002340826712),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.000396583046, - 0.002349708046),
    to_complex(0.009416709999, - 0.001604209999),
    to_complex(0.000405541339, 0.002358666339),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.000414577764, - 0.002367702764),
    to_complex(0.009489002604, - 0.001676502604),
    to_complex(0.000423693523, 0.002376818523),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.000432889836, - 0.002386014836),
    to_complex(0.009562574363, - 0.001750074363),
    to_complex(0.000442167954, 0.002395292954),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.000451529149, - 0.002404654149),
    to_complex(0.009637465219, - 0.001824965219),
    to_complex(0.000460974720, 0.002414099720),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.000470505993, - 0.002423630993),
    to_complex(0.009713716762, - 0.001901216762),
    to_complex(0.000480124323, 0.002433249323),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.000489831091, - 0.002442956091),
    to_complex(0.009791372317, - 0.001978872317),
    to_complex(0.000499627708, 0.002452752708),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.000509515614, - 0.002462640614),
    to_complex(0.009870477034, - 0.002057977034),
    to_complex(0.000519496279, 0.002472621279),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.000529571207, - 0.002482696207),
    to_complex(0.009951077986, - 0.002138577986),
    to_complex(0.000539741930, 0.002492866930),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.000550010015, - 0.002503135015),
    to_complex(0.010033224273, - 0.002220724273),
    to_complex(0.000560377065, 0.002513502065),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.000570844714, - 0.002523969714),
    to_complex(0.010116967136, - 0.002304467136),
    to_complex(0.000581414634, 0.002534539634),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.000592088532, - 0.002545213532),
    to_complex(0.010202360070, - 0.002389860070),
    to_complex(0.000602868155, 0.002555993155),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.000613755288, - 0.002566880288),
    to_complex(0.010289458953, - 0.002476958953),
    to_complex(0.000624751754, 0.002577876754),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.000635859419, - 0.002588984419),
    to_complex(0.010378322181, - 0.002565822181),
    to_complex(0.000647080190, 0.002600205190),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.000658416020, - 0.002611541020),
    to_complex(0.010469010811, - 0.002656510811),
    to_complex(0.000669868902, 0.002622993902),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.000681440879, - 0.002634565879),
    to_complex(0.010561588717, - 0.002749088717),
    to_complex(0.000693134040, 0.002646259040),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.000704950520, - 0.002658075520),
    to_complex(0.010656122748, - 0.002843622748),
    to_complex(0.000716892508, 0.002670017508),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.000728962243, - 0.002682087243),
    to_complex(0.010752682915, - 0.002940182915),
    to_complex(0.000741162015, 0.002694287015),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.000753494172, - 0.002706619172),
    to_complex(0.010851342571, - 0.003038842571),
    to_complex(0.000765961115, 0.002719086115),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.000778565306, - 0.002731690306),
    to_complex(0.010952178618, - 0.003139678618),
    to_complex(0.000791309265, 0.002744434265),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.000804195572, - 0.002757320572),
    to_complex(0.011055271724, - 0.003242771724),
    to_complex(0.000817226874, 0.002770351874),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.000830405881, - 0.002783530881),
    to_complex(0.011160706556, - 0.003348206556),
    to_complex(0.000843735370, 0.002796860370),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.000857218190, - 0.002810343190),
    to_complex(0.011268572034, - 0.003456072034),
    to_complex(0.000870857260, 0.002823982260),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.000884655572, - 0.002837780572),
    to_complex(0.011378961600, - 0.003566461600),
    to_complex(0.000898616196, 0.002851741196),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.000912742281, - 0.002865867281),
    to_complex(0.011491973509, - 0.003679473509),
    to_complex(0.000927037056, 0.002880162056),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.000941503836, - 0.002894628836),
    to_complex(0.011607711147, - 0.003795211147),
    to_complex(0.000956146021, 0.002909271021),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.000970967100, - 0.002924092100),
    to_complex(0.011726283367, - 0.003913783367),
    to_complex(0.000985970658, 0.002939095658),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.001001160372, - 0.002954285372),
    to_complex(0.011847804858, - 0.004035304858),
    to_complex(0.001016540021, 0.002969665021),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.001032113483, - 0.002985238483),
    to_complex(0.011972396542, - 0.004159896542),
    to_complex(0.001047884745, 0.003001009745),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.001063857902, - 0.003016982902),
    to_complex(0.012100186005, - 0.004287686005),
    to_complex(0.001080037162, 0.003033162162),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.001096426850, - 0.003049551850),
    to_complex(0.012231307960, - 0.004418807960),
    to_complex(0.001113031414, 0.003066156414),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.001129855426, - 0.003082980426),
    to_complex(0.012365904754, - 0.004553404754),
    to_complex(0.001146903587, 0.003100028587),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.001164180736, - 0.003117305736),
    to_complex(0.012504126920, - 0.004691626920),
    to_complex(0.001181691848, 0.003134816848),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.001199442046, - 0.003152567046),
    to_complex(0.012646133770, - 0.004833633770),
    to_complex(0.001217436599, 0.003170561599),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.001235680936, - 0.003188805936),
    to_complex(0.012792094048, - 0.004979594048),
    to_complex(0.001254180643, 0.003207305643),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.001272941476, - 0.003226066476),
    to_complex(0.012942186641, - 0.005129686641),
    to_complex(0.001291969363, 0.003245094363),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.001311270415, - 0.003264395415),
    to_complex(0.013096601347, - 0.005284101347),
    to_complex(0.001330850926, 0.003283975926),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.001350717387, - 0.003303842387),
    to_complex(0.013255539729, - 0.005443039729),
    to_complex(0.001370876491, 0.003324001491),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.001391335139, - 0.003344460139),
    to_complex(0.013419216035, - 0.005606716035),
    to_complex(0.001412100452, 0.003365225452),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.001433179777, - 0.003386304777),
    to_complex(0.013587858215, - 0.005775358215),
    to_complex(0.001454580696, 0.003407705696),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.001476311039, - 0.003429436039),
    to_complex(0.013761709038, - 0.005949209038),
    to_complex(0.001498378888, 0.003451503888),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.001520792594, - 0.003473917594),
    to_complex(0.013941027311, - 0.006128527311),
    to_complex(0.001543560783, 0.003496685783),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.001566692372, - 0.003519817372),
    to_complex(0.014126089233, - 0.006313589233),
    to_complex(0.001590196575, 0.003543321575),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.001614082923, - 0.003567207923),
    to_complex(0.014317189876, - 0.006504689876),
    to_complex(0.001638361273, 0.003591486273),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.001663041823, - 0.003616166823),
    to_complex(0.014514644829, - 0.006702144829),
    to_complex(0.001688135127, 0.003641260127),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.001713652112, - 0.003666777112),
    to_complex(0.014718792015, - 0.006906292015),
    to_complex(0.001739604090, 0.003692729090),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.001766002783, - 0.003719127783),
    to_complex(0.014929993699, - 0.007117493699),
    to_complex(0.001792860334, 0.003745985334),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.001820189331, - 0.003773314331),
    to_complex(0.015148638727, - 0.007336138727),
    to_complex(0.001848002826, 0.003801127826),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.001876314355, - 0.003829439355),
    to_complex(0.015375145004, - 0.007562645004),
    to_complex(0.001905137964, 0.003858262964),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.001934488230, - 0.003887613230),
    to_complex(0.015609962267, - 0.007797462267),
    to_complex(0.001964380289, 0.003917505289),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.001994829860, - 0.003947954860),
    to_complex(0.015853575171, - 0.008041075171),
    to_complex(0.002025853278, 0.003978978278),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.002057467519, - 0.004010592519),
    to_complex(0.016106506750, - 0.008294006750),
    to_complex(0.002089690236, 0.004042815236),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.002122539791, - 0.004075664791),
    to_complex(0.016369322293, - 0.008556822293),
    to_complex(0.002156035291, 0.004109160291),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.002190196627, - 0.004143321627),
    to_complex(0.016642633696, - 0.008830133696),
    to_complex(0.002225044515, 0.004178169515),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.002260600538, - 0.004213725538),
    to_complex(0.016927104375, - 0.009114604375),
    to_complex(0.002296887193, 0.004250012193),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.002333927938, - 0.004287052938),
    to_complex(0.017223454802, - 0.009410954802),
    to_complex(0.002371747245, 0.004324872245),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.002410370658, - 0.004363495658),
    to_complex(0.017532468773, - 0.009719968773),
    to_complex(0.002449824848, 0.004402949848),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.002490137678, - 0.004443262678),
    to_complex(0.017855000528, - 0.010042500528),
    to_complex(0.002531338269, 0.004484463269),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.002573457077, - 0.004526582077),
    to_complex(0.018191982843, - 0.010379482843),
    to_complex(0.002616525961, 0.004569650961),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.002660578275, - 0.004613703275),
    to_complex(0.018544436275, - 0.010731936275),
    to_complex(0.002705648947, 0.004658773947),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.002751774583, - 0.004704899583),
    to_complex(0.018913479732, - 0.011100979732),
    to_complex(0.002798993560, 0.004752118560),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.002847346139, - 0.004800471139),
    to_complex(0.019300342622, - 0.011487842622),
    to_complex(0.002896874583, 0.004849999583),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.002947623279, - 0.004900748279),
    to_complex(0.019706378832, - 0.011893878832),
    to_complex(0.002999638878, 0.004952763878),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.003052970435, - 0.005006095435),
    to_complex(0.020133082903, - 0.012320582903),
    to_complex(0.003107669574, 0.005060794574),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.003163790650, - 0.005116915650),
    to_complex(0.020582108778, - 0.012769608778),
    to_complex(0.003221390940, 0.005174515940),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.003280530834, - 0.005233655834),
    to_complex(0.021055291641, - 0.013242791641),
    to_complex(0.003341274056, 0.005294399056),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.003403687895, - 0.005356812895),
    to_complex(0.021554673440, - 0.013742173440),
    to_complex(0.003467843456, 0.005420968456),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.003533815938, - 0.005486940938),
    to_complex(0.022082532858, - 0.014270032858),
    to_complex(0.003601684928, 0.005554809928),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.003671534732, - 0.005624659732),
    to_complex(0.022641420645, - 0.014828920645),
    to_complex(0.003743454726, 0.005696579726),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.003817539744, - 0.005770664744),
    to_complex(0.023234201470, - 0.015421701470),
    to_complex(0.003893890499, 0.005847015499),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.003972614051, - 0.005925739051),
    to_complex(0.023864103757, - 0.016051603757),
    to_complex(0.004053824308, 0.006006949308),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.004137642590, - 0.006090767590),
    to_complex(0.024534779311, - 0.016722279311),
    to_complex(0.004224198236, 0.006177323236),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.004313629280, - 0.006266754280),
    to_complex(0.025250375081, - 0.017437875081),
    to_complex(0.004406083193, 0.006359208193),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.004501717707, - 0.006454842707),
    to_complex(0.026015620025, - 0.018203120025),
    to_complex(0.004600701718, 0.006553826718),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.004703216296, - 0.006656341296),
    to_complex(0.026835930933, - 0.019023430933),
    to_complex(0.004809455801, 0.006762580801),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.004919629121, - 0.006872754121),
    to_complex(0.027717542202, - 0.019905042202),
    to_complex(0.005033961062, 0.006987086062),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.005152693889, - 0.007105818889),
    to_complex(0.028667666156, - 0.020855166156),
    to_complex(0.005276089058, 0.007229214058),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.005404429149, - 0.007357554149),
    to_complex(0.029694692621, - 0.021882192621),
    to_complex(0.005538020051, 0.007491145051),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.005677193408, - 0.007630318408),
    to_complex(0.030808439456, - 0.022995939456),
    to_complex(0.005822309394, 0.007775434394),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.005973759849, - 0.007926884849),
    to_complex(0.032020469896, - 0.024207969896),
    to_complex(0.006131971829, 0.008085096829),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.006297411662, - 0.008250536662),
    to_complex(0.033344498452, - 0.025531998452),
    to_complex(0.006470589566, 0.008423714566),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.006652064936, - 0.008605189936),
    to_complex(0.034796915612, - 0.026984415612),
    to_complex(0.006842452413, 0.008795577413),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.007042428882, - 0.008995553882),
    to_complex(0.036397473994, - 0.028584973994),
    to_complex(0.007252741554, 0.009205866554),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.007474217340, - 0.009427342340),
    to_complex(0.038170197021, - 0.030357697021),
    to_complex(0.007707773773, 0.009660898773),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.007954431767, - 0.009907556767),
    to_complex(0.040144599158, - 0.032332099158),
    to_complex(0.008215330605, 0.010168455605),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.008491745603, - 0.010444870603),
    to_complex(0.042357349863, - 0.034544849863),
    to_complex(0.008785109036, 0.010738234036),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.009097035057, - 0.011050160057),
    to_complex(0.044854581647, - 0.037042081647),
    to_complex(0.009429349511, 0.011382474511),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.009784125813, - 0.011737250813),
    to_complex(0.047695153199, - 0.039882653199),
    to_complex(0.010163728385, 0.012116853385),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.010570865562, - 0.012523990562),
    to_complex(0.050955362780, - 0.043142862780),
    to_complex(0.011008654486, 0.012961779486),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.011480701260, - 0.013433826260),
    to_complex(0.054735924060, - 0.046923424060),
    to_complex(0.011991200739, 0.013944325739),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.012545061796, - 0.014498186796),
    to_complex(0.059172581505, - 0.051360081505),
    to_complex(0.013148065990, 0.015101190990),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.013807070518, - 0.015760195518),
    to_complex(0.064452791713, - 0.056640291713),
    to_complex(0.014530270569, 0.016483395569),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.015327542393, - 0.017280667393),
    to_complex(0.070842940328, - 0.063030440328),
    to_complex(0.016210897645, 0.018164022645),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.017195093499, - 0.019148218499),
    to_complex(0.078734770882, - 0.070922270882),
    to_complex(0.018298464629, 0.020251589629),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.019544077231, - 0.021497202231),
    to_complex(0.088728956729, - 0.080916456729),
    to_complex(0.020961360594, 0.022914485594),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.022588463793, - 0.024541588793),
    to_complex(0.101795816292, - 0.093983316292),
    to_complex(0.024475743603, 0.026428868603),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.026691072202, - 0.028644197202),
    to_complex(0.119611354027, - 0.111798854027),
    to_complex(0.029328177833, 0.031281302833),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.032520253260, - 0.034473378260),
    to_complex(0.145341356024, - 0.137528856024),
    to_complex(0.036463170193, 0.038416295193),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.041457265253, - 0.043410390253),
    to_complex(0.185769649482, - 0.177957149482),
    to_complex(0.047987697593, 0.049940822593),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.056892469387, - 0.058845594387),
    to_complex(0.258534184926, - 0.250721684926),
    to_complex(0.069754473622, 0.071707598622),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.089965623841, - 0.091918748841),
    to_complex(0.428307447286, - 0.420494947286),
    to_complex(0.126344895250, 0.128298020250),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.211228530259, - 0.213181655259),
    to_complex(1.277141799991, - 1.269329299991),
    to_complex(0.635642710525, 0.637595835525));

  -----------------------------------------------------------------------------------------------------
  constant INPUT_DATA_2048_16QAM_NOISY : complex_array(0 to 2047) := (
    to_complex(0.030235423497, - 0.057346819888),
    to_complex(- 0.003271854839, - 0.016833211267),
    to_complex(0.013845156779, 0.022982216655),
    to_complex(- 0.021945030290, - 0.037052777542),
    to_complex(- 0.024605826087, - 0.016354169205),
    to_complex(0.023345969246, 0.080726128396),
    to_complex(0.039275746679, - 0.030217787933),
    to_complex(0.068647478640, - 0.050922483932),
    to_complex(0.075462791125, - 0.002061533066),
    to_complex(- 0.045280170830, - 0.026371613966),
    to_complex(0.012696297394, 0.019282701110),
    to_complex(- 0.024791314970, - 0.015052912189),
    to_complex(- 0.060951284695, - 0.081488418409),
    to_complex(0.084219393668, 0.052933508746),
    to_complex(- 0.001591267747, - 0.053658992750),
    to_complex(- 0.004504184246, - 0.045918110289),
    to_complex(0.005007559331, 0.035892287444),
    to_complex(- 0.011091173459, - 0.041190181219),
    to_complex(0.022278954520, 0.027211831336),
    to_complex(0.026324425265, - 0.067982187418),
    to_complex(- 0.065542414419, - 0.021395217226),
    to_complex(0.078691346469, 0.138975146429),
    to_complex(- 0.000119343495, 0.009273446071),
    to_complex(0.073715369518, 0.003138313445),
    to_complex(0.052144692310, 0.082611845226),
    to_complex(- 0.017542969296, 0.039324696681),
    to_complex(- 0.002103044601, - 0.036348990591),
    to_complex(- 0.062268002700, 0.080629337981),
    to_complex(0.034509218535, - 0.021270545991),
    to_complex(0.128876019332, - 0.036827168727),
    to_complex(- 0.030419543934, - 0.063274821088),
    to_complex(0.030766453766, 0.052612561115),
    to_complex(0.097396049881, 0.050400321614),
    to_complex(0.058544813671, - 0.089844137302),
    to_complex(0.023166103829, - 0.000463741437),
    to_complex(0.000257041332, 0.027785458285),
    to_complex(- 0.010597174006, - 0.067345442271),
    to_complex(- 0.019536777763, - 0.042696996550),
    to_complex(- 0.085251995447, - 0.005501949916),
    to_complex(- 0.001618202080, - 0.074297374906),
    to_complex(0.063788917288, 0.048988039213),
    to_complex(0.085020684589, 0.035312257489),
    to_complex(0.015776687195, - 0.008376621416),
    to_complex(0.115796926063, 0.050222124882),
    to_complex(- 0.049687168420, 0.000619276571),
    to_complex(0.000439313720, - 0.030583182378),
    to_complex(0.088359022678, - 0.006804961005),
    to_complex(0.058764502294, - 0.054710249106),
    to_complex(0.035785561205, 0.001861693329),
    to_complex(- 0.014770921516, - 0.012440058569),
    to_complex(- 0.073184284357, - 0.042232297476),
    to_complex(- 0.019433941644, 0.038886066498),
    to_complex(0.027184260271, - 0.020381305718),
    to_complex(0.061508673830, 0.060114275814),
    to_complex(- 0.036704073598, 0.014183657165),
    to_complex(- 0.115533035970, - 0.095163755516),
    to_complex(- 0.017717222687, - 0.042527434415),
    to_complex(0.013805204298, - 0.012361335825),
    to_complex(0.030622082248, - 0.011913600602),
    to_complex(0.028881599340, - 0.060589813896),
    to_complex(- 0.068840147019, 0.069504010928),
    to_complex(0.021824423062, 0.122431319717),
    to_complex(- 0.027818898729, 0.067322164396),
    to_complex(- 0.024879974147, - 0.014700225655),
    to_complex(0.097480147600, - 0.001743342153),
    to_complex(0.037033634395, 0.019610797309),
    to_complex(0.023053152929, - 0.040914039839),
    to_complex(- 0.052523061125, - 0.016156587895),
    to_complex(0.076169760239, - 0.092926615426),
    to_complex(- 0.048662472433, - 0.030405420628),
    to_complex(0.034124470427, 0.008987028177),
    to_complex(- 0.009247303964, 0.017404039335),
    to_complex(0.052501469704, - 0.039503863278),
    to_complex(0.021298240218, - 0.054017647586),
    to_complex(- 0.021570784036, 0.007031604049),
    to_complex(- 0.069486287111, - 0.064848265722),
    to_complex(- 0.007060093819, 0.083537665149),
    to_complex(0.007478763853, - 0.059041893561),
    to_complex(0.063110309275, - 0.005107904445),
    to_complex(- 0.013158943439, - 0.059115290187),
    to_complex(0.041488756897, - 0.029277974512),
    to_complex(0.064314052509, - 0.036511524270),
    to_complex(- 0.036916676269, 0.054739930593),
    to_complex(- 0.059180345130, 0.023463637032),
    to_complex(- 0.057103483627, - 0.058523738175),
    to_complex(0.019806805034, 0.039112957383),
    to_complex(- 0.024700032424, - 0.074916981226),
    to_complex(- 0.000428306262, - 0.013920523280),
    to_complex(- 0.093504141067, - 0.024159668699),
    to_complex(0.065348758131, - 0.092894659896),
    to_complex(0.043765475256, - 0.024743539562),
    to_complex(- 0.047148168107, - 0.058644180881),
    to_complex(0.038002322704, - 0.031082906714),
    to_complex(0.019981466925, - 0.034502024952),
    to_complex(0.033490053342, 0.043006913453),
    to_complex(0.053790261138, 0.028695403412),
    to_complex(0.013738789399, - 0.018524956514),
    to_complex(- 0.086274650368, 0.024169151605),
    to_complex(0.048829822056, - 0.020219681460),
    to_complex(0.046178214916, - 0.103823402116),
    to_complex(0.014051969616, 0.102387483202),
    to_complex(0.031268418047, 0.078523966336),
    to_complex(0.017287682222, 0.065992001870),
    to_complex(- 0.023874620994, 0.071158568806),
    to_complex(- 0.012522581972, - 0.072377564869),
    to_complex(0.003254458085, - 0.026989914035),
    to_complex(- 0.035126768951, 0.089731760676),
    to_complex(0.050921153414, 0.084910349758),
    to_complex(- 0.029573510204, 0.005953634209),
    to_complex(- 0.006728372430, 0.030847229762),
    to_complex(- 0.095899172602, - 0.076889852282),
    to_complex(0.044561297919, - 0.100470313730),
    to_complex(- 0.019757063728, - 0.034814980847),
    to_complex(- 0.001887049047, 0.020067239344),
    to_complex(- 0.046782027552, - 0.061656611445),
    to_complex(- 0.004171651614, 0.089078836972),
    to_complex(0.027062433960, 0.036855076685),
    to_complex(0.044789551285, 0.004924986332),
    to_complex(- 0.053154069482, - 0.035411697968),
    to_complex(- 0.000337770268, 0.030938909702),
    to_complex(- 0.061994090200, 0.043657184471),
    to_complex(0.024851429897, 0.088046070585),
    to_complex(0.026380095853, - 0.019602379665),
    to_complex(- 0.029856163443, - 0.056457517966),
    to_complex(0.023978586857, - 0.022240583033),
    to_complex(0.014551043303, 0.056840729935),
    to_complex(- 0.065524514103, - 0.107193907934),
    to_complex(- 0.037836122067, 0.070431462779),
    to_complex(0.074990186432, - 0.079340374559),
    to_complex(0.077801980457, 0.008831021656),
    to_complex(- 0.026178896836, 0.034911248068),
    to_complex(- 0.021988537896, - 0.060695736047),
    to_complex(0.038957790380, 0.004944417051),
    to_complex(0.058343259388, - 0.027495149280),
    to_complex(0.062468431879, 0.040448477378),
    to_complex(- 0.054828738527, - 0.045723840993),
    to_complex(- 0.035289914240, 0.028836492399),
    to_complex(- 0.038735795547, - 0.078662478026),
    to_complex(0.057986651277, 0.039130893900),
    to_complex(- 0.085417876052, 0.024097716609),
    to_complex(- 0.058789320171, - 0.004488415239),
    to_complex(- 0.074891516937, - 0.030416935628),
    to_complex(- 0.030185925703, 0.012893114980),
    to_complex(- 0.018271667521, - 0.036573589924),
    to_complex(- 0.067046282560, 0.004420608214),
    to_complex(0.027047592993, - 0.025608414953),
    to_complex(- 0.001383778766, 0.041233581002),
    to_complex(- 0.074843567656, - 0.033436705931),
    to_complex(- 0.047371104377, - 0.001634474732),
    to_complex(0.001679938933, - 0.090980592248),
    to_complex(0.007720293805, - 0.023553372619),
    to_complex(- 0.009434425975, 0.054772569283),
    to_complex(0.064200974225, - 0.022416151112),
    to_complex(- 0.011186667921, - 0.043721303462),
    to_complex(- 0.053487548817, 0.040904301949),
    to_complex(- 0.020402018125, - 0.065607582190),
    to_complex(0.080128982654, - 0.055877507261),
    to_complex(0.065514191676, - 0.016026657873),
    to_complex(0.018420141089, - 0.010976814712),
    to_complex(0.067175030800, - 0.049860656296),
    to_complex(0.015791336437, 0.016293938271),
    to_complex(0.043167159346, - 0.007776256067),
    to_complex(0.031245212417, - 0.019941367186),
    to_complex(0.033611789890, - 0.085135835124),
    to_complex(- 0.022960351175, - 0.007953264113),
    to_complex(- 0.012046237590, 0.030200126401),
    to_complex(- 0.016772252619, - 0.065232715433),
    to_complex(0.093786397481, - 0.011386918347),
    to_complex(0.005405325314, - 0.073920486887),
    to_complex(- 0.009906781614, - 0.054831127922),
    to_complex(- 0.081904555663, 0.030705411783),
    to_complex(- 0.041046422635, 0.056355944197),
    to_complex(0.109241510608, - 0.010985169824),
    to_complex(0.029141929673, 0.048260137920),
    to_complex(0.009905040156, - 0.031785246625),
    to_complex(0.094156182455, - 0.077618409969),
    to_complex(0.069932345832, 0.074009059339),
    to_complex(0.020699036392, 0.037777385258),
    to_complex(- 0.000629819280, 0.055241622715),
    to_complex(0.031331436917, - 0.007300711311),
    to_complex(- 0.004238224933, 0.013048392564),
    to_complex(- 0.048156103508, 0.081939945780),
    to_complex(- 0.050294984401, - 0.044139884222),
    to_complex(- 0.091105700210, - 0.083512529219),
    to_complex(0.005882962085, - 0.008370316200),
    to_complex(- 0.012840616282, 0.026479196853),
    to_complex(- 0.057175276892, - 0.080029553884),
    to_complex(0.053194987711, - 0.038999593110),
    to_complex(- 0.004185746487, 0.127193130046),
    to_complex(- 0.068841710651, - 0.033919501377),
    to_complex(0.001546649295, - 0.057578163859),
    to_complex(- 0.086763826462, - 0.165632163523),
    to_complex(- 0.052390033845, 0.064321233435),
    to_complex(- 0.024032729740, - 0.028132783434),
    to_complex(0.107643118311, 0.075840324141),
    to_complex(- 0.026558032685, 0.015528193368),
    to_complex(0.054716742810, 0.078848278019),
    to_complex(0.028079390826, - 0.033406164018),
    to_complex(0.011426077114, 0.090757511562),
    to_complex(- 0.056370768160, - 0.003757789317),
    to_complex(0.053679647744, - 0.029077273660),
    to_complex(0.025698708161, 0.013014314773),
    to_complex(- 0.050081199637, 0.015645558621),
    to_complex(0.018001390053, 0.019269673595),
    to_complex(0.008695862362, 0.059869370545),
    to_complex(- 0.086626225185, - 0.032440200766),
    to_complex(0.038509216020, 0.066816409831),
    to_complex(- 0.065611286513, - 0.030013107089),
    to_complex(0.037346169060, 0.063732484161),
    to_complex(0.005846223328, 0.108487902482),
    to_complex(0.070500765945, - 0.047164148783),
    to_complex(- 0.021979565934, 0.016169584824),
    to_complex(- 0.000122480387, - 0.047807752814),
    to_complex(0.043033158552, 0.007807761125),
    to_complex(- 0.038197124507, - 0.080643482568),
    to_complex(0.136496102354, - 0.002037607528),
    to_complex(- 0.064024645180, 0.016231424177),
    to_complex(- 0.028044271404, - 0.013750851650),
    to_complex(0.080065865229, - 0.039834424272),
    to_complex(0.087877792124, - 0.046515954705),
    to_complex(- 0.009183944086, - 0.056183077437),
    to_complex(0.033921780001, - 0.017608987514),
    to_complex(- 0.056433204435, - 0.050263664959),
    to_complex(- 0.026653013316, - 0.054185533644),
    to_complex(- 0.004185072022, - 0.026965027404),
    to_complex(0.020118946053, - 0.044289813442),
    to_complex(- 0.033065357485, 0.011974699998),
    to_complex(0.090015848305, - 0.009981554838),
    to_complex(0.021197311482, - 0.030838156650),
    to_complex(0.016182706082, 0.048254451235),
    to_complex(- 0.033467788945, - 0.100633100866),
    to_complex(- 0.016718183493, 0.111893822214),
    to_complex(0.023081548988, - 0.062517268868),
    to_complex(0.042044611710, 0.082236970235),
    to_complex(0.096511202886, 0.008129680947),
    to_complex(0.004736042255, - 0.015572081794),
    to_complex(- 0.092225553543, 0.033377383841),
    to_complex(0.058240085882, - 0.050619617436),
    to_complex(0.046386543502, - 0.047209006116),
    to_complex(0.032711152912, 0.045070278157),
    to_complex(- 0.025498076138, - 0.005744206660),
    to_complex(0.015618127618, 0.035266728633),
    to_complex(0.037548222558, - 0.042624249179),
    to_complex(- 0.024491419978, - 0.045263914784),
    to_complex(0.010709496783, 0.027338205174),
    to_complex(- 0.067174815818, - 0.056998752596),
    to_complex(- 0.002313710700, 0.135659838092),
    to_complex(0.005817967858, - 0.069552726983),
    to_complex(0.056766227885, 0.024193006836),
    to_complex(0.083575300791, 0.060902339073),
    to_complex(0.025148951512, - 0.008600546558),
    to_complex(- 0.024694540918, 0.122807548153),
    to_complex(0.011488260031, - 0.025072192995),
    to_complex(- 0.016117570184, - 0.125922669694),
    to_complex(- 0.001862281002, 0.020000164405),
    to_complex(0.021244609632, 0.057294091063),
    to_complex(0.034063084847, 0.060061031076),
    to_complex(0.053854299861, 0.004443307562),
    to_complex(0.045972933705, - 0.019808711351),
    to_complex(0.090909081924, - 0.006236952645),
    to_complex(0.083384705720, 0.002225597184),
    to_complex(- 0.020736008705, - 0.067939791549),
    to_complex(- 0.024572183340, 0.020899857523),
    to_complex(- 0.029814590597, - 0.006463669604),
    to_complex(- 0.096121866079, - 0.038656587723),
    to_complex(0.023547523081, - 0.050492339236),
    to_complex(- 0.048903856773, - 0.012792738068),
    to_complex(- 0.019174675338, - 0.088727306281),
    to_complex(0.041219334780, 0.096046601515),
    to_complex(0.048092161405, 0.016157702271),
    to_complex(0.010601765777, 0.043332269517),
    to_complex(- 0.106976075365, - 0.032144484157),
    to_complex(0.034527880409, 0.072474876222),
    to_complex(- 0.088272174224, - 0.020858442563),
    to_complex(- 0.062792811240, - 0.092902642320),
    to_complex(- 0.096198781245, - 0.006095156640),
    to_complex(- 0.093147478167, - 0.056237662903),
    to_complex(0.015259263299, 0.085962428497),
    to_complex(0.103708133264, - 0.081010514105),
    to_complex(0.019535228514, 0.002580334501),
    to_complex(- 0.034282989188, - 0.006170283010),
    to_complex(0.025282369537, - 0.018430104256),
    to_complex(0.010662577103, - 0.000080542505),
    to_complex(0.190094036642, 0.012321068141),
    to_complex(- 0.022221493643, 0.011570491437),
    to_complex(0.116791519424, 0.141421796769),
    to_complex(- 0.022892591465, 0.006755744864),
    to_complex(0.020482324998, 0.040210141209),
    to_complex(- 0.022788570245, - 0.089925461734),
    to_complex(0.099812047844, 0.017342807058),
    to_complex(- 0.003069413736, 0.110447801602),
    to_complex(0.087118886463, 0.028090752631),
    to_complex(0.030764077921, - 0.015826445783),
    to_complex(0.002141864213, - 0.003413424179),
    to_complex(0.018892011944, - 0.028238539737),
    to_complex(0.034897784109, 0.036012864694),
    to_complex(0.006963074890, - 0.008592835913),
    to_complex(- 0.057226543270, - 0.014847121707),
    to_complex(- 0.027447902417, 0.026829593488),
    to_complex(0.012378314965, - 0.089783771136),
    to_complex(0.059148312753, 0.086637597633),
    to_complex(0.009248173110, 0.028179832787),
    to_complex(- 0.022268474296, 0.039909897433),
    to_complex(0.025584958447, 0.051394310621),
    to_complex(0.018398864637, 0.001233665178),
    to_complex(0.049690288937, 0.028682977244),
    to_complex(- 0.052742813016, - 0.000949138647),
    to_complex(0.060209646852, - 0.038976917155),
    to_complex(- 0.018607484818, 0.067735640313),
    to_complex(- 0.031710008124, - 0.037858624469),
    to_complex(0.017413133904, - 0.038569159665),
    to_complex(- 0.008250314998, - 0.024098554412),
    to_complex(0.006745663754, 0.047232324027),
    to_complex(0.022664957689, - 0.083646888471),
    to_complex(0.023587981503, 0.020411299513),
    to_complex(0.037817493348, - 0.026400709857),
    to_complex(0.065924583413, 0.041205498453),
    to_complex(- 0.061978069453, 0.006152533101),
    to_complex(- 0.004110001804, - 0.071023141155),
    to_complex(0.016569296153, 0.020048057568),
    to_complex(0.059321595636, - 0.031487617988),
    to_complex(- 0.037551119718, - 0.004163169994),
    to_complex(- 0.059291925359, 0.003209030036),
    to_complex(- 0.010200178013, 0.033931055927),
    to_complex(- 0.068599117695, - 0.024662056113),
    to_complex(0.012468322631, 0.091781454959),
    to_complex(0.038378886885, - 0.017162672207),
    to_complex(0.070971599040, - 0.005923518845),
    to_complex(0.065754622449, - 0.034310661818),
    to_complex(- 0.027875151498, 0.027520856083),
    to_complex(- 0.050845038193, - 0.019483902471),
    to_complex(0.078135961972, 0.053959117747),
    to_complex(- 0.063427223939, 0.065515387391),
    to_complex(0.083815724134, - 0.021380544946),
    to_complex(- 0.007711033402, 0.076156321560),
    to_complex(0.098020332706, - 0.080576105856),
    to_complex(- 0.048426868544, 0.011147015879),
    to_complex(- 0.082507695092, 0.043893421729),
    to_complex(0.011533706427, 0.002820276427),
    to_complex(- 0.077503390451, - 0.015785437747),
    to_complex(- 0.030731156491, - 0.028033194602),
    to_complex(- 0.021656895688, - 0.003782187520),
    to_complex(- 0.074994996658, - 0.024102784708),
    to_complex(0.070101412341, - 0.023450330530),
    to_complex(- 0.041128413170, - 0.075004285150),
    to_complex(- 0.051356306482, - 0.021677725999),
    to_complex(- 0.055659427012, 0.018272177544),
    to_complex(- 0.074801619351, 0.095826350502),
    to_complex(0.066344880384, 0.071936331273),
    to_complex(- 0.035202593551, 0.051086270600),
    to_complex(0.015865515739, - 0.000651192010),
    to_complex(- 0.009339754735, 0.003170348222),
    to_complex(0.029138139438, 0.061660235251),
    to_complex(- 0.001161191005, 0.007678809233),
    to_complex(0.039925864991, - 0.016067080406),
    to_complex(- 0.016187873507, 0.054962878043),
    to_complex(- 0.042001828267, - 0.060140666784),
    to_complex(0.004789074013, 0.058201574131),
    to_complex(- 0.096439779457, 0.090066039720),
    to_complex(0.055368445662, - 0.066047181942),
    to_complex(0.092543579393, - 0.021938448646),
    to_complex(0.041262164040, - 0.024883579374),
    to_complex(0.002224827122, - 0.067799453359),
    to_complex(- 0.023043571970, 0.091144162957),
    to_complex(- 0.062325795597, - 0.033286912218),
    to_complex(0.026751297060, 0.097003952378),
    to_complex(- 0.050461860392, - 0.020295778445),
    to_complex(- 0.004583565271, 0.049064994918),
    to_complex(- 0.068247273024, - 0.134821711276),
    to_complex(0.015708878116, 0.055245620757),
    to_complex(0.038977418417, 0.012676655629),
    to_complex(- 0.001836268521, - 0.014629410047),
    to_complex(- 0.031435003133, 0.016813534030),
    to_complex(- 0.082305899838, 0.001503603851),
    to_complex(- 0.030317498894, 0.142886575418),
    to_complex(0.070366673001, 0.019243692286),
    to_complex(- 0.029982253756, 0.073554346322),
    to_complex(- 0.049350079722, 0.063949244570),
    to_complex(- 0.031213558752, 0.045050266132),
    to_complex(0.058103536764, 0.021634948193),
    to_complex(0.042081864891, - 0.036313003747),
    to_complex(- 0.019920774686, 0.054566579998),
    to_complex(- 0.051337740308, - 0.050465385685),
    to_complex(0.010570220042, 0.004725926254),
    to_complex(- 0.105674606224, 0.016387342440),
    to_complex(- 0.014947853373, 0.068781008606),
    to_complex(0.019128243796, 0.023643299160),
    to_complex(- 0.120016241544, 0.058419057738),
    to_complex(0.006791687635, 0.024023821022),
    to_complex(- 0.030113640872, - 0.013211846017),
    to_complex(0.078466063974, - 0.050023866972),
    to_complex(0.058479564103, - 0.077723783065),
    to_complex(- 0.025959360791, - 0.044491530958),
    to_complex(0.031218323935, - 0.038539717809),
    to_complex(0.117937831000, - 0.005580457443),
    to_complex(0.041713003278, - 0.018605568589),
    to_complex(0.027161156988, - 0.015963227212),
    to_complex(0.036071145463, - 0.015303213708),
    to_complex(- 0.036917798255, - 0.052644290896),
    to_complex(0.109769640844, 0.017789337162),
    to_complex(0.045166482693, 0.064237596497),
    to_complex(- 0.024353791653, - 0.063258782882),
    to_complex(- 0.033762453902, - 0.027378687709),
    to_complex(0.001563122782, 0.138856686658),
    to_complex(0.007670442611, - 0.057263058562),
    to_complex(- 0.053082416674, 0.018628316578),
    to_complex(0.007732009257, 0.139237473695),
    to_complex(0.000043997191, 0.032481162821),
    to_complex(0.032726379958, - 0.026850263142),
    to_complex(- 0.073752106138, 0.000510084538),
    to_complex(- 0.048527428012, 0.062529344123),
    to_complex(- 0.147297258296, 0.006456423121),
    to_complex(0.087310399464, - 0.011380516914),
    to_complex(- 0.000390464533, - 0.098592454821),
    to_complex(0.028690182836, - 0.034797348894),
    to_complex(- 0.049950792763, - 0.104292752993),
    to_complex(- 0.057748691874, 0.057847309970),
    to_complex(0.000795643649, 0.025296250801),
    to_complex(0.082059795320, - 0.005510954094),
    to_complex(0.050879542563, - 0.009365642652),
    to_complex(0.034101416516, - 0.003568086166),
    to_complex(- 0.039865513674, 0.034410208972),
    to_complex(0.029077070486, 0.000677339422),
    to_complex(0.044652182246, - 0.009280387865),
    to_complex(0.022616096462, 0.033834694768),
    to_complex(0.038148122232, - 0.097891797922),
    to_complex(0.051469949409, - 0.018424327254),
    to_complex(- 0.052160890892, 0.032478272383),
    to_complex(- 0.052403996265, - 0.034002607438),
    to_complex(- 0.037371978827, - 0.037388403863),
    to_complex(0.101893428275, - 0.132617171163),
    to_complex(- 0.021860310324, 0.034115403360),
    to_complex(0.001044937131, - 0.060233959532),
    to_complex(- 0.021385069551, 0.058645727125),
    to_complex(- 0.075219264605, - 0.051854005253),
    to_complex(0.001400793052, 0.061026621375),
    to_complex(- 0.013563439464, - 0.047357052366),
    to_complex(- 0.003721054293, 0.011363335816),
    to_complex(0.034413771233, - 0.083220242222),
    to_complex(0.015267682121, - 0.036055165206),
    to_complex(0.051235399666, - 0.024671870586),
    to_complex(0.086742297623, - 0.012814850862),
    to_complex(0.027357983043, - 0.018947979154),
    to_complex(- 0.018808547113, 0.028156294716),
    to_complex(0.029321251911, - 0.057549655592),
    to_complex(- 0.004604189498, 0.049299380902),
    to_complex(- 0.000707299578, 0.014516355199),
    to_complex(0.018442453083, - 0.003657022960),
    to_complex(0.069901258990, 0.020296960641),
    to_complex(0.052796870257, 0.055059308083),
    to_complex(- 0.005498587975, - 0.086537864676),
    to_complex(- 0.023183579673, - 0.014040750207),
    to_complex(- 0.120284498995, - 0.091818964265),
    to_complex(- 0.026690635160, - 0.044427342640),
    to_complex(- 0.043612681472, 0.049345461857),
    to_complex(- 0.026444212283, - 0.083309804583),
    to_complex(- 0.032660966977, 0.016121711055),
    to_complex(0.028200254379, - 0.000982353231),
    to_complex(0.029667540265, 0.013240901107),
    to_complex(0.076927881279, 0.015536431666),
    to_complex(- 0.032117894932, - 0.043048629251),
    to_complex(- 0.022233462276, 0.035254605293),
    to_complex(0.101593399168, 0.068284011517),
    to_complex(- 0.063444148586, - 0.078529460702),
    to_complex(0.029722013268, - 0.024458302982),
    to_complex(0.008708134422, 0.078987207976),
    to_complex(- 0.035146365175, 0.008248874543),
    to_complex(0.031041965442, - 0.037629476567),
    to_complex(- 0.131029337615, - 0.057737965003),
    to_complex(- 0.016002677966, - 0.043625591979),
    to_complex(0.039598255756, 0.036941584312),
    to_complex(0.024289240422, 0.067460206057),
    to_complex(- 0.020264214243, - 0.085522282442),
    to_complex(0.099719064091, 0.045791719747),
    to_complex(0.105743110047, - 0.008943893497),
    to_complex(0.044174002834, 0.087335840220),
    to_complex(- 0.020010232998, - 0.035652184208),
    to_complex(0.044366221689, - 0.010629623337),
    to_complex(- 0.122625768797, 0.019990546058),
    to_complex(0.063108964224, 0.012098572770),
    to_complex(0.035895196017, 0.004690424614),
    to_complex(- 0.025877027440, - 0.010185223561),
    to_complex(- 0.000887638464, 0.032391866051),
    to_complex(0.064935026404, - 0.072089797018),
    to_complex(- 0.008898318960, - 0.049547705538),
    to_complex(- 0.057072769188, 0.016838555590),
    to_complex(0.051088304536, - 0.077086510345),
    to_complex(- 0.071240958004, - 0.006332196341),
    to_complex(0.036909249163, - 0.109109663560),
    to_complex(- 0.067264943800, - 0.061765208137),
    to_complex(- 0.057234056963, - 0.002076278595),
    to_complex(- 0.020323252996, 0.027491094463),
    to_complex(0.013648619796, - 0.065004084073),
    to_complex(0.046437168944, 0.014246972140),
    to_complex(0.044687138012, 0.023554152532),
    to_complex(- 0.023134733348, 0.055615611555),
    to_complex(- 0.072662886159, - 0.010316666051),
    to_complex(- 0.006975915411, - 0.040783526943),
    to_complex(- 0.000173228852, 0.032418596483),
    to_complex(- 0.009221239516, 0.004175239458),
    to_complex(- 0.045006873675, - 0.049108901715),
    to_complex(0.027557086152, 0.013645816036),
    to_complex(- 0.013823443583, 0.053124721816),
    to_complex(0.025943494433, - 0.034780689319),
    to_complex(- 0.041457148804, 0.044497357901),
    to_complex(- 0.003171857478, 0.020321732980),
    to_complex(- 0.050799332330, - 0.043545372526),
    to_complex(0.049525447305, - 0.075491983187),
    to_complex(- 0.072887060759, - 0.107635062828),
    to_complex(- 0.039916142258, - 0.079219860199),
    to_complex(- 0.018871310309, - 0.020627554399),
    to_complex(- 0.025909736744, 0.056126832534),
    to_complex(0.079451118245, 0.006489967271),
    to_complex(0.020764215229, - 0.026528468535),
    to_complex(- 0.005319220985, - 0.069216497344),
    to_complex(- 0.000244175339, 0.009354627908),
    to_complex(- 0.002176592368, 0.021824298350),
    to_complex(- 0.048637432737, - 0.031445299754),
    to_complex(- 0.005300932586, - 0.039874479514),
    to_complex(0.046346052606, - 0.060237550797),
    to_complex(0.034860527200, - 0.057436977111),
    to_complex(0.112963131496, - 0.044885819579),
    to_complex(0.050640656659, - 0.026347018736),
    to_complex(- 0.040123149331, - 0.035374042595),
    to_complex(0.013831719168, - 0.010540726244),
    to_complex(0.069345245909, 0.049802440153),
    to_complex(0.008997888173, - 0.024207516891),
    to_complex(0.002604685858, 0.069397731223),
    to_complex(- 0.017995568718, - 0.039478346913),
    to_complex(0.042281840196, 0.015262407812),
    to_complex(0.007240819216, - 0.041301946394),
    to_complex(0.046556615491, 0.046539175697),
    to_complex(0.020830404412, 0.095779292949),
    to_complex(0.029387463374, 0.019353451127),
    to_complex(- 0.000220758808, 0.056845624847),
    to_complex(0.064981314597, - 0.010347440311),
    to_complex(- 0.039076494226, - 0.153831269422),
    to_complex(0.024535594286, - 0.027513938210),
    to_complex(0.047771954863, 0.021363940892),
    to_complex(0.033863470822, 0.056157316418),
    to_complex(- 0.121168348040, - 0.004677922635),
    to_complex(- 0.074910435898, - 0.040498943643),
    to_complex(- 0.088908427722, 0.066271567498),
    to_complex(- 0.006126896171, - 0.034591511464),
    to_complex(0.048925816426, - 0.008847704585),
    to_complex(0.043841334119, 0.003533842028),
    to_complex(0.063106192275, - 0.026167711284),
    to_complex(- 0.021275329941, - 0.045069599501),
    to_complex(0.009856207527, - 0.006010403059),
    to_complex(0.050883588301, - 0.009461287253),
    to_complex(- 0.025886865619, 0.021000374860),
    to_complex(0.077432531843, - 0.121067547720),
    to_complex(0.004419050172, - 0.094577743109),
    to_complex(0.088298377032, 0.008397487377),
    to_complex(0.049658027953, 0.018839453367),
    to_complex(0.044057176679, - 0.032227256832),
    to_complex(- 0.025268248598, 0.020636349504),
    to_complex(- 0.043279112626, 0.094342075977),
    to_complex(- 0.030083435414, - 0.101473356151),
    to_complex(- 0.031718695854, - 0.028188360640),
    to_complex(0.071367204482, 0.014908269420),
    to_complex(0.083217238395, 0.024043834771),
    to_complex(0.027914412051, 0.012650182139),
    to_complex(- 0.058568473080, 0.030280193907),
    to_complex(0.028435863196, - 0.066867283353),
    to_complex(0.029774368383, - 0.034950165170),
    to_complex(0.083440026473, - 0.022024044296),
    to_complex(- 0.011857254186, 0.062428604571),
    to_complex(- 0.121646922103, 0.021985587055),
    to_complex(- 0.113897814357, 0.073672084448),
    to_complex(0.027373441201, 0.040110233916),
    to_complex(0.007752036367, 0.004465961924),
    to_complex(0.007501282105, 0.014881027925),
    to_complex(- 0.026400878439, 0.045209006411),
    to_complex(- 0.061138893436, 0.006407088851),
    to_complex(0.002072741376, 0.089141692567),
    to_complex(- 0.028915481049, 0.055514324660),
    to_complex(0.049777772576, 0.055826720235),
    to_complex(0.042544481578, 0.032735327126),
    to_complex(0.068365378696, 0.024482889711),
    to_complex(- 0.009920819917, 0.023538067089),
    to_complex(0.021338928115, 0.000126610168),
    to_complex(- 0.004673397729, 0.007140468226),
    to_complex(0.002361246250, - 0.015393323101),
    to_complex(0.035265889147, 0.049218027806),
    to_complex(0.093272738882, 0.030368246011),
    to_complex(- 0.021671253965, 0.018044644784),
    to_complex(- 0.092686863740, - 0.001371657294),
    to_complex(- 0.038762245701, 0.003520714402),
    to_complex(- 0.034787322191, 0.018789446782),
    to_complex(- 0.012516142474, - 0.022465385762),
    to_complex(0.057672350595, 0.072927257823),
    to_complex(- 0.048255178843, - 0.023966498371),
    to_complex(0.079442561890, - 0.017484062970),
    to_complex(- 0.020129667283, - 0.112482077319),
    to_complex(- 0.060471183017, - 0.023744956026),
    to_complex(0.035026704890, - 0.010727397975),
    to_complex(- 0.016365732298, - 0.061275452899),
    to_complex(- 0.072028652410, 0.000461414924),
    to_complex(0.092109558907, - 0.002067901930),
    to_complex(- 0.024774803435, 0.069667644311),
    to_complex(0.039821365067, 0.050194282829),
    to_complex(- 0.049245461127, - 0.014679107648),
    to_complex(0.010929036370, 0.015644936498),
    to_complex(0.019599272149, 0.044414403853),
    to_complex(- 0.061705537701, 0.034621484734),
    to_complex(- 0.047762487549, - 0.042008900502),
    to_complex(- 0.046022936283, - 0.027736951501),
    to_complex(- 0.025466813163, 0.028634585491),
    to_complex(- 0.013629294972, - 0.045567711856),
    to_complex(0.006418825946, 0.049441163281),
    to_complex(0.012271517593, - 0.077651018689),
    to_complex(0.094757126208, - 0.024568684756),
    to_complex(- 0.000569246136, - 0.012144488450),
    to_complex(0.098465907674, - 0.084613519883),
    to_complex(- 0.036732929870, - 0.006849256178),
    to_complex(- 0.001543440229, 0.016584175376),
    to_complex(0.026515493422, - 0.037275589129),
    to_complex(0.031710139791, 0.047206559975),
    to_complex(0.146187488861, 0.009739884488),
    to_complex(- 0.058736939820, - 0.073525643758),
    to_complex(0.024505565854, - 0.002482063604),
    to_complex(- 0.074681162234, 0.005841436252),
    to_complex(- 0.065378742172, 0.035079425854),
    to_complex(- 0.057007950295, - 0.012659051440),
    to_complex(0.054086353233, - 0.002550317805),
    to_complex(0.034698957026, - 0.014473244856),
    to_complex(- 0.010319634742, 0.014416668631),
    to_complex(- 0.005442103345, 0.059675176067),
    to_complex(- 0.007371305196, - 0.009337347357),
    to_complex(- 0.051544440839, - 0.011554306489),
    to_complex(0.074558065836, 0.014511209586),
    to_complex(- 0.094894029873, 0.001037952721),
    to_complex(0.073029537938, - 0.062628992774),
    to_complex(0.075703909305, 0.051855337822),
    to_complex(0.050699777189, - 0.031252696464),
    to_complex(- 0.019478568248, - 0.019311962539),
    to_complex(- 0.044561903266, - 0.040488278929),
    to_complex(0.074642964100, 0.057409482648),
    to_complex(0.059537751798, - 0.107646633655),
    to_complex(- 0.057274493801, 0.119546961245),
    to_complex(- 0.057253101214, 0.028192206226),
    to_complex(0.040846551353, 0.041407307098),
    to_complex(0.040848268143, 0.007574125082),
    to_complex(0.013168821849, 0.042663861175),
    to_complex(- 0.029058858479, - 0.022394761159),
    to_complex(0.017652016375, 0.001664658495),
    to_complex(- 0.006120968967, 0.018487981584),
    to_complex(0.062596759295, - 0.006090436381),
    to_complex(- 0.055682514941, 0.027113005750),
    to_complex(0.042085127662, - 0.037535479221),
    to_complex(- 0.054465328782, 0.005331356467),
    to_complex(0.003235395726, - 0.077134526241),
    to_complex(- 0.013587287321, - 0.055662275728),
    to_complex(- 0.046461086877, 0.052051959696),
    to_complex(- 0.018929539380, - 0.053866624439),
    to_complex(- 0.001393942732, - 0.016226766107),
    to_complex(0.021488721873, - 0.037683867977),
    to_complex(0.039010978690, 0.021342334429),
    to_complex(0.057038271381, 0.017136971378),
    to_complex(- 0.043225335804, 0.099909155421),
    to_complex(0.006497204422, 0.018883276115),
    to_complex(- 0.093259861068, - 0.011327787958),
    to_complex(- 0.015937355156, 0.111946916937),
    to_complex(0.010310876727, - 0.057362670355),
    to_complex(0.013050477116, - 0.038086440142),
    to_complex(- 0.059825628980, 0.040644472848),
    to_complex(- 0.003792567829, 0.026387693507),
    to_complex(0.066496619173, 0.009500376975),
    to_complex(0.054145813274, - 0.016964317625),
    to_complex(- 0.076422289378, 0.025690019278),
    to_complex(- 0.012975063429, - 0.033359516108),
    to_complex(0.006564283756, 0.012407606313),
    to_complex(- 0.045700068092, - 0.001914531768),
    to_complex(- 0.019903982404, - 0.095601984489),
    to_complex(- 0.054332410012, - 0.051073660261),
    to_complex(- 0.009864436383, 0.003576062492),
    to_complex(- 0.098421532237, 0.107475708791),
    to_complex(- 0.018145733200, - 0.041124251864),
    to_complex(0.088321562061, 0.103277462930),
    to_complex(- 0.051847140888, - 0.040030695263),
    to_complex(0.066965566052, 0.010944725220),
    to_complex(- 0.020033957482, 0.086916019984),
    to_complex(0.019372572002, 0.046439147432),
    to_complex(- 0.024410325932, - 0.011857088624),
    to_complex(- 0.009279557043, 0.004313548213),
    to_complex(- 0.036220964686, - 0.014796587542),
    to_complex(0.043415439391, - 0.017532628716),
    to_complex(0.049034242107, 0.002903457408),
    to_complex(0.049805062655, 0.095732426109),
    to_complex(- 0.052375495997, - 0.017858021345),
    to_complex(- 0.063584740540, - 0.013366685865),
    to_complex(- 0.019333774576, - 0.011316514745),
    to_complex(0.001923717741, - 0.011932537865),
    to_complex(- 0.000649999089, 0.010835256297),
    to_complex(- 0.106841414531, 0.004070270769),
    to_complex(- 0.061190917478, - 0.080406888760),
    to_complex(0.056742376663, - 0.013600221985),
    to_complex(- 0.010593258449, 0.041676589130),
    to_complex(- 0.050182932408, - 0.057367548770),
    to_complex(0.050482012461, - 0.043906268706),
    to_complex(- 0.062873235001, 0.015823789058),
    to_complex(0.043422788757, - 0.101128411969),
    to_complex(0.033480624000, - 0.050935743449),
    to_complex(- 0.015987629653, 0.007852391772),
    to_complex(- 0.093872714620, 0.001783444062),
    to_complex(- 0.015460508226, - 0.027124108728),
    to_complex(- 0.066021360911, - 0.074337084338),
    to_complex(0.051962600562, 0.106189789055),
    to_complex(0.045360631581, 0.057155357702),
    to_complex(- 0.048110154132, - 0.055131808150),
    to_complex(- 0.053132084787, 0.070631939301),
    to_complex(- 0.056046143331, - 0.046657038822),
    to_complex(0.080306999890, 0.074742868829),
    to_complex(0.051460674087, 0.048673832729),
    to_complex(0.060638090914, 0.030874754799),
    to_complex(- 0.004544872201, 0.031148150171),
    to_complex(0.048482726355, 0.024062169416),
    to_complex(- 0.037479085121, - 0.006930644462),
    to_complex(- 0.027862910545, 0.078257352958),
    to_complex(- 0.108446458166, 0.093836788837),
    to_complex(0.023074241280, - 0.002992166283),
    to_complex(0.065702987683, - 0.002058222280),
    to_complex(- 0.017093211398, 0.026273894402),
    to_complex(- 0.063872573185, 0.022862172948),
    to_complex(0.008118257959, - 0.031158107851),
    to_complex(- 0.005959794630, - 0.013323421570),
    to_complex(- 0.063194649043, - 0.027321896792),
    to_complex(- 0.025730131620, 0.014947352719),
    to_complex(0.046211269848, - 0.002685082104),
    to_complex(- 0.018788794913, 0.048130191020),
    to_complex(0.051962309380, 0.017424211168),
    to_complex(- 0.071004791576, 0.078893983658),
    to_complex(- 0.006343466574, - 0.046044948334),
    to_complex(- 0.027928954070, 0.083814586923),
    to_complex(0.042933890373, - 0.061704891172),
    to_complex(0.034477936694, - 0.068220770162),
    to_complex(- 0.002025509363, 0.018667167781),
    to_complex(0.011023672066, - 0.030359581313),
    to_complex(- 0.035696285349, 0.033839615088),
    to_complex(0.053124509259, 0.039843131387),
    to_complex(0.005379880112, 0.016156748924),
    to_complex(- 0.095982227027, - 0.031628058440),
    to_complex(0.017637431875, - 0.002891621861),
    to_complex(0.072860626685, 0.036307544247),
    to_complex(- 0.012790366338, 0.019209228065),
    to_complex(- 0.066589341692, - 0.010454853115),
    to_complex(0.011984821667, 0.123123396896),
    to_complex(0.042866093896, 0.096804601219),
    to_complex(- 0.020996338964, 0.026895641109),
    to_complex(- 0.043764685108, 0.016145960805),
    to_complex(0.005453201844, 0.011225153567),
    to_complex(- 0.003494555190, - 0.022145524925),
    to_complex(- 0.013714201639, - 0.024247372986),
    to_complex(0.000963574622, - 0.032826832400),
    to_complex(- 0.003989409163, - 0.067110231301),
    to_complex(- 0.032490713142, 0.031092534328),
    to_complex(- 0.114424500242, - 0.009733281571),
    to_complex(- 0.014108019981, 0.045056477375),
    to_complex(0.068246946306, 0.052539561751),
    to_complex(- 0.068552598957, - 0.013225447615),
    to_complex(0.017128115750, 0.097743982613),
    to_complex(- 0.027664419625, - 0.068499708160),
    to_complex(- 0.040482797178, 0.073203254277),
    to_complex(0.010384401041, 0.119827333996),
    to_complex(0.023064492781, 0.035740909701),
    to_complex(- 0.025279563323, - 0.039862612434),
    to_complex(- 0.033082925539, 0.056927150722),
    to_complex(0.086423015296, 0.068000107559),
    to_complex(0.011160790247, 0.039804375217),
    to_complex(- 0.028196002163, 0.059436115849),
    to_complex(0.025434523765, 0.096090022472),
    to_complex(0.061108533889, 0.013801208057),
    to_complex(- 0.029830800003, 0.022268386603),
    to_complex(0.029726139286, 0.021321575390),
    to_complex(- 0.041070582864, - 0.031506680564),
    to_complex(- 0.021149966300, - 0.044115357228),
    to_complex(0.008927542384, 0.053278253621),
    to_complex(- 0.008409639377, - 0.013497112882),
    to_complex(- 0.002010076219, - 0.035213141788),
    to_complex(0.021474115041, 0.064303728609),
    to_complex(0.013686824923, 0.001023296133),
    to_complex(- 0.055575507091, 0.077442527405),
    to_complex(0.052868766100, 0.035739198439),
    to_complex(- 0.013677910384, - 0.041763414586),
    to_complex(0.033285500053, 0.018259209371),
    to_complex(- 0.024931404842, - 0.052058481655),
    to_complex(0.095579295718, - 0.035519723414),
    to_complex(- 0.087477652136, - 0.056579746554),
    to_complex(- 0.025876479123, 0.054278552327),
    to_complex(- 0.023325430920, 0.095784938194),
    to_complex(- 0.065768132081, 0.086570711669),
    to_complex(0.061464012596, - 0.060599601699),
    to_complex(0.019538453682, - 0.013940823167),
    to_complex(0.038049601853, - 0.013321729376),
    to_complex(- 0.080541023913, 0.002921235923),
    to_complex(0.013025027240, - 0.058385407375),
    to_complex(- 0.019654101389, 0.040016235833),
    to_complex(- 0.025851434315, - 0.023119192476),
    to_complex(- 0.010915493475, - 0.022956710929),
    to_complex(0.083440727902, 0.030822358322),
    to_complex(0.069921307619, - 0.045409766743),
    to_complex(- 0.006567350372, - 0.052837120906),
    to_complex(- 0.009943865355, - 0.033007999603),
    to_complex(- 0.069620335234, - 0.099844678325),
    to_complex(- 0.084849267316, - 0.048962287108),
    to_complex(- 0.030350998087, 0.041156890308),
    to_complex(- 0.070910409682, - 0.025617734651),
    to_complex(0.032687919443, - 0.007900037336),
    to_complex(0.058753048801, - 0.006535435178),
    to_complex(0.025350946209, - 0.039872171444),
    to_complex(- 0.040680013146, 0.010824136656),
    to_complex(0.056811991493, 0.023706110783),
    to_complex(- 0.003331034292, 0.080891738241),
    to_complex(0.047210687375, - 0.026383006000),
    to_complex(- 0.029334275193, - 0.003141160276),
    to_complex(- 0.015503253802, 0.053818733081),
    to_complex(0.009650201409, - 0.001471711372),
    to_complex(- 0.075521100993, 0.020984632770),
    to_complex(0.038952025287, 0.027233106234),
    to_complex(- 0.056959245475, 0.031950170006),
    to_complex(- 0.107810189929, - 0.019153288750),
    to_complex(0.073619943372, - 0.087940186330),
    to_complex(0.072818295537, 0.011656535948),
    to_complex(- 0.048688573729, - 0.024354513580),
    to_complex(- 0.010504908762, 0.046722749105),
    to_complex(- 0.004756525349, 0.051665945923),
    to_complex(- 0.062700376677, - 0.035384151086),
    to_complex(0.067787306293, - 0.014758050728),
    to_complex(- 0.014801659663, - 0.013096353766),
    to_complex(- 0.002631336649, 0.045322300080),
    to_complex(0.033747885857, 0.032594927894),
    to_complex(0.055715444577, 0.136345536978),
    to_complex(0.071479494509, 0.002069717962),
    to_complex(- 0.011744619421, - 0.014131846575),
    to_complex(- 0.049028096783, 0.043133211507),
    to_complex(- 0.078078285555, 0.013260624306),
    to_complex(0.043125548220, - 0.035659021924),
    to_complex(0.002966108879, 0.036849037055),
    to_complex(- 0.089589334093, 0.019429636084),
    to_complex(0.020718159814, - 0.014694754737),
    to_complex(0.045470996853, - 0.043992557408),
    to_complex(- 0.015116683674, - 0.107979716588),
    to_complex(- 0.003928318998, 0.003941247218),
    to_complex(- 0.029069657876, - 0.068886012439),
    to_complex(- 0.018221809704, 0.051145102624),
    to_complex(0.026813357272, - 0.053044443678),
    to_complex(0.067227449997, 0.062009063716),
    to_complex(- 0.002365591143, 0.040707948118),
    to_complex(0.037036968781, - 0.035976151714),
    to_complex(0.002523521625, - 0.076623309179),
    to_complex(0.008334168984, - 0.022325658320),
    to_complex(- 0.063696163287, - 0.048942820141),
    to_complex(0.013161066436, - 0.073837902136),
    to_complex(- 0.076439426840, 0.004516373407),
    to_complex(0.039273451441, 0.040248880237),
    to_complex(- 0.023814438623, - 0.020446522049),
    to_complex(0.095022395282, 0.016920168314),
    to_complex(- 0.096836497751, - 0.005725244013),
    to_complex(0.051005050761, 0.017454394823),
    to_complex(- 0.035551685388, - 0.028938112200),
    to_complex(0.035223557708, - 0.005553488163),
    to_complex(0.037156683257, 0.003868590226),
    to_complex(- 0.001732307140, 0.054574377160),
    to_complex(- 0.012535589947, - 0.031691473404),
    to_complex(0.051214717373, 0.021186732938),
    to_complex(- 0.053930378486, - 0.002664012843),
    to_complex(0.013986184699, - 0.035884075216),
    to_complex(- 0.019484149943, - 0.014550314514),
    to_complex(0.031585363603, - 0.063314240498),
    to_complex(0.063956675125, - 0.065376090093),
    to_complex(- 0.011494152871, 0.016033841149),
    to_complex(- 0.038587082865, - 0.005926039416),
    to_complex(0.047527146941, 0.137416757255),
    to_complex(0.022051707072, - 0.059536228535),
    to_complex(- 0.069198984684, 0.034278995048),
    to_complex(0.031846568089, - 0.014444846771),
    to_complex(- 0.039092025498, - 0.008088694512),
    to_complex(- 0.027776795968, - 0.014062476158),
    to_complex(0.068389460425, 0.106325242145),
    to_complex(0.002943752653, - 0.013297274805),
    to_complex(0.018144380927, 0.067041839791),
    to_complex(- 0.042853457149, - 0.009103198678),
    to_complex(- 0.016429808852, 0.054338823049),
    to_complex(- 0.150853688494, 0.029266910748),
    to_complex(0.040809179197, - 0.018181853968),
    to_complex(0.105132537631, 0.049192310738),
    to_complex(0.007515220512, 0.037567676359),
    to_complex(0.085254615331, - 0.011972828961),
    to_complex(- 0.067640228122, - 0.010133212417),
    to_complex(0.103842628418, 0.022718709559),
    to_complex(0.186306150038, - 0.053895405544),
    to_complex(0.088854609765, 0.084497005145),
    to_complex(- 0.061829371775, 0.055277895969),
    to_complex(- 0.014621177146, 0.044848107589),
    to_complex(- 0.004477237284, - 0.093069727104),
    to_complex(- 0.027919811400, - 0.056814331027),
    to_complex(- 0.063363613194, - 0.107474350631),
    to_complex(- 0.040005020853, 0.031403781622),
    to_complex(0.039331882727, 0.010656099296),
    to_complex(- 0.000176872037, 0.003476481253),
    to_complex(- 0.053630808702, 0.010047244874),
    to_complex(- 0.130779750193, 0.060086941304),
    to_complex(- 0.009066657615, - 0.009188103942),
    to_complex(0.045803540259, 0.055244495757),
    to_complex(- 0.031783294646, 0.005940837908),
    to_complex(0.014057720008, - 0.004110936134),
    to_complex(- 0.044701870093, 0.039052925647),
    to_complex(- 0.001391237855, - 0.045862360526),
    to_complex(- 0.026360545067, - 0.019278697486),
    to_complex(0.019898282966, 0.035417263625),
    to_complex(- 0.011100324846, - 0.062706030981),
    to_complex(0.003356253073, - 0.006677011600),
    to_complex(- 0.030486919780, - 0.040241965704),
    to_complex(0.000916324431, - 0.037769877353),
    to_complex(0.055854730304, 0.030946939459),
    to_complex(- 0.052519738465, - 0.041504864343),
    to_complex(- 0.016863186684, 0.014595500974),
    to_complex(0.020809826397, - 0.015409219474),
    to_complex(0.071534187747, 0.012383780863),
    to_complex(0.004047596486, 0.020500854004),
    to_complex(0.027939033800, 0.078043006241),
    to_complex(- 0.011186207261, 0.031463965721),
    to_complex(- 0.061030511962, - 0.061829681379),
    to_complex(- 0.102883684092, 0.070220697463),
    to_complex(- 0.125854741604, 0.013695288410),
    to_complex(- 0.087159409109, - 0.036390191696),
    to_complex(- 0.003138745619, 0.028831032244),
    to_complex(0.002519853174, - 0.024797453225),
    to_complex(- 0.033361256087, 0.058304860468),
    to_complex(- 0.037325571019, - 0.074011215043),
    to_complex(- 0.005339982691, 0.081747727700),
    to_complex(0.025515022503, - 0.027172586714),
    to_complex(- 0.038163187138, - 0.006942772109),
    to_complex(0.025840481245, 0.037842869981),
    to_complex(0.074451684307, 0.073076463563),
    to_complex(- 0.001209552900, 0.045714903570),
    to_complex(0.017601982509, - 0.013067003350),
    to_complex(- 0.089355479995, 0.043921192255),
    to_complex(0.066472844008, - 0.032678649660),
    to_complex(- 0.056886062088, 0.020708040584),
    to_complex(- 0.024198124153, 0.017632695854),
    to_complex(0.013478716126, - 0.054545362680),
    to_complex(0.089861096260, - 0.015191390586),
    to_complex(- 0.001970160065, 0.077362850019),
    to_complex(- 0.021881561542, 0.040138742689),
    to_complex(0.012348974419, - 0.045168288583),
    to_complex(0.082242017144, 0.027551893595),
    to_complex(- 0.039192418798, - 0.059051747373),
    to_complex(- 0.042027829218, 0.048867558277),
    to_complex(0.047016104970, - 0.071067940698),
    to_complex(0.000774909076, 0.099612584228),
    to_complex(- 0.009606022576, - 0.058124045166),
    to_complex(0.034422891611, 0.011448513966),
    to_complex(- 0.010482158309, - 0.075778519313),
    to_complex(- 0.028667817338, 0.042303443508),
    to_complex(0.021073769676, - 0.008537239478),
    to_complex(0.065502392686, - 0.056491315305),
    to_complex(0.036721511025, 0.065663005658),
    to_complex(0.078588679811, - 0.001015165291),
    to_complex(0.055445603711, - 0.011191337208),
    to_complex(- 0.057020889584, - 0.014904918546),
    to_complex(- 0.029859426061, 0.024650522946),
    to_complex(- 0.083996535580, - 0.009993678546),
    to_complex(- 0.013937228000, - 0.031900063210),
    to_complex(- 0.042832308919, 0.005720774063),
    to_complex(0.017674314034, - 0.050687565008),
    to_complex(0.012548582956, 0.025344253023),
    to_complex(- 0.020457905163, 0.007418060672),
    to_complex(0.034142903473, - 0.002980277491),
    to_complex(- 0.014631383573, 0.031591067156),
    to_complex(- 0.054291442521, 0.019965655408),
    to_complex(- 0.132360908069, - 0.020720230755),
    to_complex(0.017618951544, - 0.003229622751),
    to_complex(- 0.028229870285, 0.000946919599),
    to_complex(- 0.020911128871, 0.072555823880),
    to_complex(- 0.066944568984, 0.027772804758),
    to_complex(0.013964075232, 0.055688624337),
    to_complex(0.011246314759, 0.009683051897),
    to_complex(- 0.010724952681, 0.053474545499),
    to_complex(- 0.007797194187, 0.004859256094),
    to_complex(- 0.017475181625, 0.056712337051),
    to_complex(0.011579851661, - 0.055721767281),
    to_complex(0.024361657072, 0.128985891550),
    to_complex(0.047127002189, 0.070383998099),
    to_complex(0.011894960903, - 0.023448114129),
    to_complex(- 0.027485161979, - 0.034145091959),
    to_complex(0.072369516899, 0.033471786443),
    to_complex(0.018280177341, 0.011757898468),
    to_complex(- 0.045803975097, 0.017422376020),
    to_complex(- 0.032443932447, 0.002772285391),
    to_complex(0.039766008944, - 0.005780652048),
    to_complex(- 0.041093244583, - 0.033250695562),
    to_complex(- 0.043827621397, - 0.014857663878),
    to_complex(- 0.034557967254, - 0.006752009936),
    to_complex(- 0.031258860273, 0.067421377492),
    to_complex(0.042305895569, - 0.002138081187),
    to_complex(0.030686091261, - 0.088483010164),
    to_complex(0.056029105653, 0.010802094888),
    to_complex(0.042026449782, 0.023487388530),
    to_complex(- 0.049941210905, 0.064419921010),
    to_complex(0.053847756296, - 0.015859404026),
    to_complex(- 0.017634904519, - 0.142095607238),
    to_complex(- 0.040473229048, 0.012953335296),
    to_complex(0.044471269653, 0.044322405402),
    to_complex(- 0.005208569196, 0.062802137100),
    to_complex(- 0.042550427468, 0.014469824262),
    to_complex(- 0.072125133233, - 0.016555620917),
    to_complex(- 0.037814672392, - 0.114018920728),
    to_complex(0.029674189540, - 0.064171474740),
    to_complex(- 0.044787537925, - 0.006201108373),
    to_complex(0.040299389462, - 0.001503936419),
    to_complex(- 0.043649452744, - 0.056047195526),
    to_complex(0.041606049928, - 0.061979997849),
    to_complex(0.025083326910, 0.023275804503),
    to_complex(- 0.070442950375, - 0.023890404923),
    to_complex(0.066804021115, - 0.050935280925),
    to_complex(0.001698684972, 0.101731310059),
    to_complex(- 0.056077552723, - 0.030626891404),
    to_complex(0.004346048332, 0.031047104386),
    to_complex(0.023964012269, - 0.041653194900),
    to_complex(0.010749419841, 0.005838970269),
    to_complex(0.024683038356, - 0.017051562422),
    to_complex(0.015135600843, - 0.073751238661),
    to_complex(- 0.019660892812, 0.026486744573),
    to_complex(0.021406587577, 0.073258681871),
    to_complex(- 0.016741075022, - 0.084210596591),
    to_complex(0.060935690277, 0.038972724224),
    to_complex(- 0.036982452908, 0.058468115481),
    to_complex(0.092220216259, - 0.021255087194),
    to_complex(0.071409159644, - 0.005295385165),
    to_complex(0.011592411277, 0.090116909836),
    to_complex(- 0.039876707483, - 0.100343396463),
    to_complex(- 0.050240048395, - 0.007465798085),
    to_complex(0.019367995602, - 0.036435332988),
    to_complex(0.077077947912, 0.064800102478),
    to_complex(0.032167618057, 0.123446894974),
    to_complex(- 0.050953909794, 0.076438358603),
    to_complex(- 0.016467663724, 0.022802201678),
    to_complex(- 0.035472226659, 0.121085082149),
    to_complex(0.027450430893, 0.057501788634),
    to_complex(- 0.086727120693, - 0.037800708863),
    to_complex(- 0.016651953887, 0.012783585319),
    to_complex(- 0.089912285951, - 0.037190353142),
    to_complex(0.026957156772, 0.046521785134),
    to_complex(- 0.014121993925, - 0.002141043490),
    to_complex(0.047735175019, - 0.013088530125),
    to_complex(- 0.070757152298, - 0.003485749405),
    to_complex(0.071790331347, 0.008251211049),
    to_complex(0.023909564352, - 0.033497914932),
    to_complex(- 0.080031164330, 0.008148796427),
    to_complex(0.048990070293, - 0.023912730509),
    to_complex(0.100828753982, 0.085980068622),
    to_complex(- 0.032545925260, 0.140719160918),
    to_complex(0.025358054228, - 0.078300131687),
    to_complex(0.022311937597, - 0.038691849878),
    to_complex(0.001802081606, 0.052201579353),
    to_complex(0.073206773472, 0.003169970017),
    to_complex(- 0.057029326016, 0.026196099267),
    to_complex(0.032134825184, 0.025576705611),
    to_complex(- 0.019886961976, 0.015533252192),
    to_complex(0.017262181347, 0.117475966951),
    to_complex(- 0.042953289826, 0.053770352149),
    to_complex(- 0.097302451971, 0.032516599353),
    to_complex(- 0.058947060136, - 0.016122832110),
    to_complex(- 0.009977132763, - 0.091078336702),
    to_complex(0.000567583546, 0.034870451150),
    to_complex(0.029397912557, - 0.020135743405),
    to_complex(- 0.029083031976, - 0.004848660811),
    to_complex(0.023818043220, - 0.105256495212),
    to_complex(0.013136464759, - 0.033182521960),
    to_complex(0.023283167287, 0.036108508673),
    to_complex(- 0.060839795188, - 0.030275175884),
    to_complex(- 0.055112593846, 0.011154750307),
    to_complex(- 0.008329090843, - 0.035907102451),
    to_complex(- 0.090478407862, - 0.053928273489),
    to_complex(0.028408417679, - 0.000156504207),
    to_complex(- 0.041874666943, 0.028314661903),
    to_complex(0.018239601637, - 0.091692039020),
    to_complex(- 0.045504346123, - 0.073956727212),
    to_complex(- 0.028998265928, 0.052332534283),
    to_complex(- 0.069588555471, - 0.003530941490),
    to_complex(0.033652186212, - 0.042125956610),
    to_complex(0.013187216724, - 0.032826099859),
    to_complex(0.066851579539, 0.021848482814),
    to_complex(- 0.016309350116, - 0.023599490603),
    to_complex(- 0.005176380597, 0.035152755295),
    to_complex(0.053404623410, - 0.057967424282),
    to_complex(0.008408108339, 0.000963213616),
    to_complex(- 0.025924391511, 0.080411414517),
    to_complex(0.042144661599, 0.012208427811),
    to_complex(0.058506267434, 0.021586985300),
    to_complex(- 0.002424941867, - 0.055849539862),
    to_complex(0.025123660854, - 0.054972347752),
    to_complex(0.058046017988, - 0.006678400581),
    to_complex(- 0.009189272336, - 0.015063813078),
    to_complex(- 0.026522983667, - 0.091387809599),
    to_complex(- 0.009182434330, 0.014084075054),
    to_complex(0.079130331366, 0.133993119118),
    to_complex(- 0.047066044753, - 0.008272209708),
    to_complex(0.034555540271, 0.138061283482),
    to_complex(- 0.084320314371, - 0.028354367940),
    to_complex(0.054001923452, 0.026191272625),
    to_complex(0.059322391577, - 0.089943321240),
    to_complex(- 0.020422401200, - 0.004447475415),
    to_complex(0.018849121771, 0.034691941978),
    to_complex(- 0.021425244655, - 0.017348439459),
    to_complex(0.046632204359, - 0.056581264294),
    to_complex(- 0.021802208524, 0.060033269704),
    to_complex(- 0.146530359167, - 0.044746490957),
    to_complex(0.099726489316, 0.004366611644),
    to_complex(0.103549320162, - 0.023581254657),
    to_complex(0.027903046305, 0.038124913993),
    to_complex(- 0.066850240606, 0.026572352897),
    to_complex(0.055393296480, 0.009314213349),
    to_complex(- 0.091199046319, - 0.004640473255),
    to_complex(- 0.002361986325, - 0.027062180184),
    to_complex(0.003821260957, 0.009839567493),
    to_complex(- 0.022217996938, 0.003571717641),
    to_complex(- 0.011479511197, - 0.015627633240),
    to_complex(0.021962447524, 0.045644907885),
    to_complex(- 0.047827991011, - 0.060729877092),
    to_complex(0.022841576410, - 0.011235632755),
    to_complex(- 0.061779243121, - 0.000877551463),
    to_complex(0.080653807424, 0.057828748963),
    to_complex(0.039505258218, 0.024913356617),
    to_complex(- 0.038135409508, - 0.001639678381),
    to_complex(0.072171604265, 0.096291976385),
    to_complex(0.073661586963, 0.010640587686),
    to_complex(0.018245464486, - 0.078174087468),
    to_complex(0.005049873748, 0.054976381277),
    to_complex(0.070660506868, - 0.058965134406),
    to_complex(- 0.015364386329, - 0.006744233624),
    to_complex(0.021411115437, 0.055305417601),
    to_complex(0.057172218060, - 0.109620659965),
    to_complex(- 0.007445944360, - 0.021341853950),
    to_complex(0.019735898280, 0.060366513321),
    to_complex(0.094575621048, - 0.003246485243),
    to_complex(- 0.022067998096, 0.032403036174),
    to_complex(- 0.018268900105, - 0.047629343262),
    to_complex(- 0.014853445873, 0.006260340026),
    to_complex(- 0.006940064890, 0.089923919024),
    to_complex(- 0.017157350434, 0.003872612724),
    to_complex(0.024036964353, - 0.063426053384),
    to_complex(0.005852064765, 0.020819995831),
    to_complex(- 0.004526893189, - 0.030558448714),
    to_complex(- 0.021882626957, 0.028530285931),
    to_complex(0.033039309210, 0.041231480023),
    to_complex(0.036103107140, - 0.033278601100),
    to_complex(0.006718168077, - 0.035169468149),
    to_complex(- 0.016109023008, - 0.067664870816),
    to_complex(0.043196031858, 0.037580666383),
    to_complex(0.006498820005, 0.074584661527),
    to_complex(- 0.082729721679, - 0.028863435079),
    to_complex(0.044273831381, 0.095166739985),
    to_complex(0.069457065213, - 0.024004257854),
    to_complex(- 0.064773419743, 0.063886629526),
    to_complex(- 0.016444541320, - 0.004023177458),
    to_complex(0.046129320815, 0.007921089842),
    to_complex(0.026982782242, 0.006328099589),
    to_complex(- 0.077404134924, 0.041592169064),
    to_complex(0.046342390272, 0.094154343264),
    to_complex(0.079477938977, 0.011720542865),
    to_complex(- 0.009632329874, - 0.166818056666),
    to_complex(- 0.043306482322, - 0.021460626329),
    to_complex(0.010177127053, - 0.022521303403),
    to_complex(- 0.015921510209, - 0.026562923725),
    to_complex(0.012108091056, 0.050875122124),
    to_complex(0.001441254219, 0.011499097016),
    to_complex(- 0.026415871339, - 0.112387879189),
    to_complex(0.020019964659, 0.021374148549),
    to_complex(0.076022045386, - 0.048573141560),
    to_complex(0.025014684440, - 0.011059506724),
    to_complex(- 0.001294944658, 0.039422829246),
    to_complex(0.008877297220, 0.054832333211),
    to_complex(- 0.006939782781, - 0.008602333591),
    to_complex(0.007890099212, 0.038054875992),
    to_complex(0.024469941583, - 0.002722362567),
    to_complex(0.007628144285, 0.045977504663),
    to_complex(- 0.016217899465, 0.012550517461),
    to_complex(- 0.052129071911, - 0.033509451316),
    to_complex(- 0.056510464689, 0.033430252668),
    to_complex(- 0.024110368304, 0.021743450632),
    to_complex(- 0.029454654444, 0.010078234515),
    to_complex(0.070504790741, - 0.007617309725),
    to_complex(- 0.099667956958, 0.009507176555),
    to_complex(- 0.001630142058, - 0.054683363153),
    to_complex(- 0.023513655006, 0.052307402655),
    to_complex(- 0.012907084527, 0.015814245641),
    to_complex(- 0.033984903860, - 0.056727616831),
    to_complex(- 0.041382189101, 0.046321019006),
    to_complex(0.056138580894, - 0.032321154757),
    to_complex(- 0.103847396323, - 0.007361584692),
    to_complex(- 0.002917896629, - 0.019452240383),
    to_complex(0.000094042649, 0.066034221619),
    to_complex(0.042523936969, - 0.085800081757),
    to_complex(0.037964778891, 0.045388513578),
    to_complex(- 0.046204638329, - 0.027728353564),
    to_complex(0.051591493828, 0.010879719277),
    to_complex(- 0.067826750522, - 0.017360354398),
    to_complex(- 0.098024273558, - 0.009255104144),
    to_complex(0.075264877424, 0.102121454671),
    to_complex(- 0.033127394964, - 0.047520804263),
    to_complex(0.007354129480, - 0.027204149691),
    to_complex(- 0.114837985468, 0.015657365564),
    to_complex(0.011553446017, 0.015599489001),
    to_complex(- 0.049803811036, 0.021162157953),
    to_complex(- 0.041095507895, 0.017116412806),
    to_complex(0.019471477707, 0.038257625726),
    to_complex(- 0.086037533382, - 0.013850644282),
    to_complex(0.084939190870, - 0.083771257809),
    to_complex(- 0.033562421922, 0.052287444256),
    to_complex(- 0.014968271836, - 0.034596749265),
    to_complex(0.066295748553, 0.044512950956),
    to_complex(- 0.085893613177, 0.007596220226),
    to_complex(0.007225889332, 0.029841747440),
    to_complex(0.001570360583, - 0.024087166426),
    to_complex(0.013889448207, - 0.026784948861),
    to_complex(0.063146025648, - 0.052920744226),
    to_complex(- 0.002772897895, 0.051273693193),
    to_complex(0.017758395632, 0.039636298025),
    to_complex(0.010134998336, 0.062599395534),
    to_complex(- 0.141944758350, 0.028853659025),
    to_complex(0.003090918259, - 0.027401753393),
    to_complex(0.087445799759, - 0.041514123516),
    to_complex(- 0.046143835146, - 0.045325732949),
    to_complex(0.022226289631, - 0.038296382898),
    to_complex(0.018630541032, 0.015062507530),
    to_complex(0.050732247872, 0.001745026589),
    to_complex(- 0.002230315508, - 0.002869656036),
    to_complex(- 0.005607448422, 0.015646343162),
    to_complex(- 0.018475402595, - 0.009107640637),
    to_complex(0.059342501605, - 0.024373094873),
    to_complex(0.041981057322, 0.109615639773),
    to_complex(- 0.057736663223, 0.053286000109),
    to_complex(0.031833521117, 0.032220113454),
    to_complex(0.054559259304, - 0.048134174969),
    to_complex(- 0.044935884431, - 0.000670544845),
    to_complex(- 0.109501219679, 0.087341443082),
    to_complex(0.056313905515, 0.018216299085),
    to_complex(- 0.038745305848, - 0.061895438706),
    to_complex(0.001219369656, 0.010466732226),
    to_complex(0.078596250997, - 0.053249117216),
    to_complex(0.093749969871, 0.006660672051),
    to_complex(0.085153104461, - 0.012994667547),
    to_complex(- 0.056245933460, 0.042712795075),
    to_complex(0.010421264801, - 0.045338704540),
    to_complex(0.040889140419, - 0.043085272704),
    to_complex(0.023076777518, 0.019912152664),
    to_complex(- 0.015907519536, - 0.014866405473),
    to_complex(- 0.084814031505, - 0.001264247819),
    to_complex(- 0.050034601583, - 0.004540585372),
    to_complex(0.055854754339, - 0.020817546857),
    to_complex(- 0.065722878872, 0.092045236286),
    to_complex(- 0.046968014639, - 0.021491452312),
    to_complex(0.010971333167, 0.073408839478),
    to_complex(0.056016272757, 0.020265792592),
    to_complex(- 0.016337183350, - 0.020800920540),
    to_complex(0.073626567474, 0.029513163237),
    to_complex(0.020430129696, - 0.078840621335),
    to_complex(- 0.108030625468, - 0.026742468783),
    to_complex(0.001984951250, - 0.043153948633),
    to_complex(0.023949628400, - 0.016629174524),
    to_complex(- 0.018730737243, - 0.023333020786),
    to_complex(- 0.068814955737, 0.036658084008),
    to_complex(- 0.052601958595, - 0.010552770087),
    to_complex(0.004222417482, - 0.003224674575),
    to_complex(0.073049215612, - 0.062141797320),
    to_complex(- 0.101611070098, - 0.005442997329),
    to_complex(- 0.036565401076, - 0.030702988266),
    to_complex(- 0.006089259622, 0.035397146441),
    to_complex(- 0.023936218886, 0.016606297764),
    to_complex(0.059872559079, 0.033919398447),
    to_complex(0.014060746578, 0.007435005920),
    to_complex(- 0.035370408485, - 0.054168065815),
    to_complex(0.021158759924, 0.002959783170),
    to_complex(- 0.072779066955, 0.084550518464),
    to_complex(0.029111532370, 0.071835407361),
    to_complex(- 0.056923839922, - 0.014349644625),
    to_complex(- 0.005640868228, - 0.054781713558),
    to_complex(- 0.021300702664, - 0.078618433753),
    to_complex(0.001619846978, 0.013172073846),
    to_complex(- 0.027154649254, 0.008094646646),
    to_complex(0.028696040646, - 0.014418459834),
    to_complex(0.021734133507, - 0.109370475355),
    to_complex(0.028253190555, - 0.012602049448),
    to_complex(- 0.070878048854, 0.072002924846),
    to_complex(- 0.051719370211, 0.008980140302),
    to_complex(0.004413233164, 0.000262664092),
    to_complex(- 0.059274292625, - 0.036424363535),
    to_complex(0.037444410752, - 0.039587313889),
    to_complex(0.018468277096, - 0.038153692389),
    to_complex(- 0.002343982232, 0.020033041370),
    to_complex(0.073919170225, - 0.047027178553),
    to_complex(- 0.030273428314, 0.024757726798),
    to_complex(0.013815344180, 0.004189961812),
    to_complex(0.000062092236, - 0.017089152413),
    to_complex(- 0.055673748932, - 0.021780549831),
    to_complex(0.058643712109, - 0.028153429048),
    to_complex(- 0.027348202415, - 0.036208142108),
    to_complex(0.004842163009, - 0.002335842026),
    to_complex(- 0.080144490993, - 0.010163850777),
    to_complex(0.028396848860, - 0.017492063879),
    to_complex(0.028747752989, 0.007810823565),
    to_complex(- 0.044374184319, - 0.039794067836),
    to_complex(0.012975207549, - 0.039889960627),
    to_complex(- 0.084672384183, 0.047401329489),
    to_complex(- 0.012762207286, 0.049462622314),
    to_complex(0.072940585690, 0.009654137180),
    to_complex(0.020680000652, 0.036348026883),
    to_complex(0.052532824649, 0.059157961350),
    to_complex(0.036487784903, 0.043427619751),
    to_complex(- 0.070357483340, - 0.033128298737),
    to_complex(- 0.006211545331, - 0.005287505316),
    to_complex(- 0.060717779118, - 0.060430752889),
    to_complex(- 0.040549800132, 0.091508781545),
    to_complex(- 0.024268510541, 0.057006266908),
    to_complex(0.025806249857, - 0.033458312805),
    to_complex(- 0.004034509236, - 0.046033381790),
    to_complex(- 0.004254795824, 0.015341586610),
    to_complex(0.089615952847, 0.058493932847),
    to_complex(- 0.092297984168, - 0.000187770081),
    to_complex(0.026287211257, 0.094693246112),
    to_complex(- 0.019194550646, - 0.019885539905),
    to_complex(- 0.053381759311, - 0.109315853588),
    to_complex(- 0.025407411519, 0.015227416002),
    to_complex(0.030237787560, 0.055132730894),
    to_complex(0.026095578741, - 0.014947644519),
    to_complex(0.013897450816, 0.066658974326),
    to_complex(0.120697642133, 0.021975591820),
    to_complex(- 0.015064015832, 0.056560741208),
    to_complex(- 0.006113556948, 0.054057401374),
    to_complex(0.028983405192, 0.005942540183),
    to_complex(0.021637817835, 0.052571590046),
    to_complex(0.028303659661, - 0.090449878784),
    to_complex(- 0.018685902349, 0.026260712100),
    to_complex(0.072823710735, - 0.014741124667),
    to_complex(0.053549610135, - 0.020912591571),
    to_complex(0.052540951255, - 0.042380918839),
    to_complex(- 0.038570406840, 0.003694470765),
    to_complex(- 0.054282261030, 0.118842451831),
    to_complex(0.031897448935, - 0.135898259248),
    to_complex(- 0.111775138662, 0.046191575899),
    to_complex(0.029403086100, 0.059812303079),
    to_complex(0.026040679642, 0.028284675319),
    to_complex(- 0.011764915368, 0.008284517290),
    to_complex(0.012175749533, 0.019964974703),
    to_complex(- 0.030825391890, 0.007262849400),
    to_complex(0.020355604281, - 0.012826750453),
    to_complex(- 0.007289028748, - 0.026767118841),
    to_complex(- 0.022807062379, 0.040001872281),
    to_complex(0.077702567703, - 0.019536571134),
    to_complex(0.030132804094, - 0.018188568555),
    to_complex(- 0.012657764435, 0.018912625734),
    to_complex(- 0.021767592584, - 0.061614107774),
    to_complex(0.047471846688, - 0.083785641405),
    to_complex(0.018448792086, 0.002668598079),
    to_complex(0.035140596843, 0.073273184353),
    to_complex(- 0.010412840317, 0.044014314208),
    to_complex(0.045661802943, - 0.016044523750),
    to_complex(0.137602655462, - 0.167619562427),
    to_complex(0.054331337543, - 0.056839403183),
    to_complex(0.059833008842, 0.062309489930),
    to_complex(0.058581171577, - 0.001470754112),
    to_complex(0.059008753229, 0.068573660554),
    to_complex(- 0.011609379784, 0.040952519865),
    to_complex(- 0.063816044834, - 0.054213806933),
    to_complex(- 0.019149250801, - 0.086315584518),
    to_complex(0.054995329706, - 0.053563026510),
    to_complex(- 0.023801057193, 0.055038706912),
    to_complex(- 0.060180372688, 0.089686855532),
    to_complex(0.031885499771, - 0.104997838319),
    to_complex(0.016732241182, 0.003962151686),
    to_complex(- 0.025815535303, 0.002273479456),
    to_complex(- 0.069123845253, 0.042410924994),
    to_complex(- 0.064510430042, - 0.001952384145),
    to_complex(0.031533593845, 0.032469688388),
    to_complex(- 0.010972483710, - 0.015853415423),
    to_complex(0.068883627836, 0.000478546083),
    to_complex(0.006422081760, - 0.040151133155),
    to_complex(- 0.020170454259, - 0.005861416828),
    to_complex(0.075937229805, - 0.012575295472),
    to_complex(- 0.006677113026, - 0.056779775191),
    to_complex(- 0.067976327436, 0.010868285581),
    to_complex(- 0.006269782125, - 0.003999257153),
    to_complex(- 0.127133910724, 0.008743958336),
    to_complex(- 0.006773271246, - 0.047464825871),
    to_complex(0.033380689732, - 0.002640565680),
    to_complex(- 0.072494459958, 0.011785716578),
    to_complex(0.055075498829, - 0.042773937782),
    to_complex(- 0.058442151142, 0.105757257422),
    to_complex(- 0.049791394025, - 0.002136700198),
    to_complex(- 0.060335855168, 0.007926026712),
    to_complex(- 0.023545829110, - 0.118675733452),
    to_complex(0.088711800169, 0.009778428148),
    to_complex(- 0.018574865723, 0.059289246804),
    to_complex(- 0.096841969458, 0.025419274160),
    to_complex(- 0.026705618149, 0.032020884930),
    to_complex(- 0.047502518043, 0.019313506660),
    to_complex(0.003920800030, - 0.054092033103),
    to_complex(- 0.026403721230, - 0.013564949654),
    to_complex(- 0.047099532166, 0.002034344200),
    to_complex(0.062029446943, - 0.000484186708),
    to_complex(0.027812500779, - 0.025496381835),
    to_complex(0.007428307950, 0.029299997297),
    to_complex(0.012319396946, - 0.036321289605),
    to_complex(0.001492830638, - 0.070944484855),
    to_complex(- 0.056251128392, - 0.079713743978),
    to_complex(0.076849363900, 0.110210927406),
    to_complex(- 0.055473655589, 0.059400683823),
    to_complex(0.066446203845, 0.013693037922),
    to_complex(- 0.068196724729, - 0.033074913562),
    to_complex(- 0.041733457509, - 0.018131486315),
    to_complex(0.007268795722, - 0.022914097703),
    to_complex(0.104545298752, 0.005085362760),
    to_complex(- 0.002608680860, - 0.048988455851),
    to_complex(0.024025477510, 0.004707069648),
    to_complex(- 0.069184499123, - 0.097452738308),
    to_complex(- 0.038897242130, 0.031029762301),
    to_complex(- 0.038082908481, - 0.026275853227),
    to_complex(0.005843382580, - 0.031984804967),
    to_complex(0.053424550909, - 0.066984593815),
    to_complex(0.018013057817, 0.038851744343),
    to_complex(0.054977036826, - 0.014110007391),
    to_complex(0.037136520403, 0.027912344906),
    to_complex(- 0.062353391957, 0.022175858370),
    to_complex(0.063785595563, 0.033657540004),
    to_complex(0.003806684463, - 0.039695460066),
    to_complex(- 0.009080697486, 0.017908186249),
    to_complex(- 0.070897299299, 0.095416153872),
    to_complex(- 0.034564500615, - 0.079584680457),
    to_complex(0.040779349054, 0.051626285974),
    to_complex(- 0.102679924418, 0.004653411767),
    to_complex(0.024432485983, - 0.019628739576),
    to_complex(- 0.066197752690, 0.115252753817),
    to_complex(0.003631104223, 0.059462279603),
    to_complex(0.038521913120, - 0.118185260300),
    to_complex(0.064341125392, 0.019891648617),
    to_complex(0.036823937205, - 0.029265662981),
    to_complex(- 0.021564055745, 0.006229004645),
    to_complex(- 0.004947153933, 0.012288018122),
    to_complex(- 0.024437603250, 0.031299117763),
    to_complex(0.109008687970, - 0.099155363728),
    to_complex(0.014595948156, - 0.074260996711),
    to_complex(0.029466018475, - 0.055557126798),
    to_complex(0.038521728606, - 0.019082877436),
    to_complex(0.049779201675, - 0.030279500790),
    to_complex(0.021158169503, - 0.095449596473),
    to_complex(0.041184813211, 0.101064168949),
    to_complex(- 0.025119911083, - 0.007006539552),
    to_complex(0.043124220140, - 0.031811842154),
    to_complex(0.040584934237, 0.038560618323),
    to_complex(0.041850488279, - 0.075412254609),
    to_complex(0.012123025249, - 0.073457390635),
    to_complex(- 0.015358075152, 0.008754551021),
    to_complex(0.030580552517, 0.055860035626),
    to_complex(0.104355449687, - 0.038307707045),
    to_complex(- 0.033394796941, - 0.066017964923),
    to_complex(0.023175844962, 0.030072336819),
    to_complex(- 0.094511540020, - 0.015254113600),
    to_complex(0.032976363177, - 0.031643431357),
    to_complex(- 0.037443488000, 0.033638435340),
    to_complex(0.016646692804, 0.002030546320),
    to_complex(- 0.066599708630, 0.089170745343),
    to_complex(- 0.077560719045, 0.042030345330),
    to_complex(0.042620058473, 0.017054664639),
    to_complex(0.078705365259, - 0.015700759350),
    to_complex(- 0.029252544542, - 0.008885907840),
    to_complex(- 0.043485542888, 0.040405812097),
    to_complex(0.074262561331, 0.042343584524),
    to_complex(- 0.047788406147, 0.058030166284),
    to_complex(0.044865403965, 0.039251620214),
    to_complex(0.006074811096, 0.003918332125),
    to_complex(- 0.014801054495, 0.011593503820),
    to_complex(- 0.001401790943, 0.008180177329),
    to_complex(0.028908962482, 0.075048513505),
    to_complex(0.006986854238, 0.063333230295),
    to_complex(- 0.014282062957, 0.024908109911),
    to_complex(0.028459420950, - 0.017016081875),
    to_complex(0.002237112422, 0.094077861717),
    to_complex(0.058343940734, 0.006957432820),
    to_complex(0.113602546846, - 0.020464998689),
    to_complex(- 0.081539767994, 0.029650993340),
    to_complex(0.034016786113, 0.008024730979),
    to_complex(- 0.048846586989, - 0.092139351418),
    to_complex(- 0.038130872772, - 0.045749145980),
    to_complex(- 0.023836258859, 0.046649857881),
    to_complex(- 0.012379656598, - 0.065529183187),
    to_complex(0.010595469521, - 0.000901595513),
    to_complex(0.058444499329, - 0.013695307451),
    to_complex(- 0.106575079556, - 0.007904846458),
    to_complex(0.042392948991, 0.055694263225),
    to_complex(0.124136909829, - 0.040731829077),
    to_complex(0.002614825808, - 0.064791922547),
    to_complex(0.037026600795, - 0.017754210404),
    to_complex(- 0.022349265307, - 0.099550605637),
    to_complex(- 0.089715279025, - 0.052170182650),
    to_complex(- 0.086162341723, - 0.053676678025),
    to_complex(- 0.074096771921, 0.049648062401),
    to_complex(0.008882317494, 0.044809081185),
    to_complex(0.017656967778, - 0.023170992712),
    to_complex(0.083789569236, - 0.021549532316),
    to_complex(0.058551954929, - 0.002304891256),
    to_complex(- 0.008913447625, 0.061968305024),
    to_complex(- 0.070153957626, 0.089755500979),
    to_complex(- 0.013368713938, 0.000811269116),
    to_complex(0.025951870049, - 0.054239772364),
    to_complex(- 0.010470737976, - 0.009074976759),
    to_complex(0.009430610242, - 0.016740962988),
    to_complex(- 0.072024063019, - 0.000036122773),
    to_complex(- 0.039908418755, - 0.043448578714),
    to_complex(0.071363904212, 0.021398175248),
    to_complex(- 0.041758652591, 0.034709906941),
    to_complex(- 0.007387292076, - 0.070833537896),
    to_complex(- 0.008118900957, - 0.024805876797),
    to_complex(- 0.033445188387, 0.038127205664),
    to_complex(0.015280630111, - 0.033147961223),
    to_complex(- 0.017848415691, - 0.008766926458),
    to_complex(- 0.011938755936, - 0.074298578719),
    to_complex(- 0.055577349079, - 0.051190640138),
    to_complex(0.062988391185, 0.071748791641),
    to_complex(- 0.017746868102, - 0.045802216890),
    to_complex(- 0.019551566190, 0.028961812139),
    to_complex(0.069332463943, - 0.083757657666),
    to_complex(0.022878283738, 0.047021402369),
    to_complex(0.028680697220, - 0.009010467863),
    to_complex(- 0.094592394152, 0.125239563031),
    to_complex(0.001783081226, 0.039628919307),
    to_complex(- 0.065852072404, 0.010348158317),
    to_complex(- 0.087137226731, 0.014920862740),
    to_complex(0.006372345077, 0.005567414293),
    to_complex(0.006795959337, - 0.022568073427),
    to_complex(0.053622285247, - 0.036392356952),
    to_complex(- 0.008178711466, - 0.057785985312),
    to_complex(0.063978508572, - 0.073377563639),
    to_complex(- 0.016014606036, 0.010702096651),
    to_complex(- 0.074341584376, - 0.028682105232),
    to_complex(0.024320703712, - 0.071835822789),
    to_complex(0.018593612425, - 0.034930119539),
    to_complex(0.030720487502, 0.071080406997),
    to_complex(0.038034923850, 0.017448509409),
    to_complex(- 0.000432064318, 0.022790510011),
    to_complex(0.065421278775, 0.007738422210),
    to_complex(- 0.062074864214, - 0.017760270755),
    to_complex(0.003423984055, - 0.040432551769),
    to_complex(0.074085941033, 0.077316672052),
    to_complex(- 0.096102129079, 0.016574028113),
    to_complex(- 0.035984555141, 0.036694977168),
    to_complex(0.021764716196, 0.042259525516),
    to_complex(0.003231100154, - 0.042798351540),
    to_complex(- 0.028253659283, 0.053354631995),
    to_complex(0.021826952281, 0.050840022653),
    to_complex(- 0.020803433877, 0.044690364262),
    to_complex(0.103478559144, 0.101188026418),
    to_complex(- 0.083221234983, 0.038004817883),
    to_complex(- 0.003634534148, - 0.025453800336),
    to_complex(0.047578267855, - 0.034326491474),
    to_complex(0.022855439438, 0.039435970965),
    to_complex(- 0.011703140568, 0.052688724289),
    to_complex(0.099025056365, 0.115737904843),
    to_complex(- 0.017846720488, - 0.065536475682),
    to_complex(- 0.042616782552, 0.121915929795),
    to_complex(0.028080647453, - 0.002146687420),
    to_complex(0.055116316406, - 0.002393303694),
    to_complex(- 0.018923872242, 0.020762569920),
    to_complex(0.006469630845, - 0.113429983574),
    to_complex(0.050660477776, 0.064011938070),
    to_complex(- 0.005662565484, - 0.001394925906),
    to_complex(- 0.009788713760, 0.038650609269),
    to_complex(0.058546269633, 0.011505357402),
    to_complex(0.003542329104, - 0.030505423470),
    to_complex(- 0.065245880687, 0.068492772703),
    to_complex(0.136848542820, - 0.022354756788),
    to_complex(0.011100466096, 0.043306369388),
    to_complex(- 0.034617457288, 0.022999358111),
    to_complex(0.041586167656, 0.068727919723),
    to_complex(0.011172902198, 0.000921303188),
    to_complex(0.054374606111, - 0.046222559949),
    to_complex(- 0.040484318560, - 0.008965187688),
    to_complex(0.037885953042, 0.024771653890),
    to_complex(0.068092956193, - 0.110185667588),
    to_complex(- 0.004421013056, - 0.053342649108),
    to_complex(- 0.009353053474, 0.018588912507),
    to_complex(0.011643596352, 0.028053445376),
    to_complex(0.056180179098, 0.074479525391),
    to_complex(- 0.029949923983, 0.093337503518),
    to_complex(- 0.061146888507, 0.106111859088),
    to_complex(0.006773000650, 0.034451792372),
    to_complex(0.020132707834, 0.025676849864),
    to_complex(- 0.040198578387, - 0.004406098586),
    to_complex(0.039794995109, 0.016853313442),
    to_complex(- 0.114398306561, 0.030969272803),
    to_complex(0.001291719673, - 0.035035768392),
    to_complex(- 0.008807617026, - 0.057804452953),
    to_complex(- 0.040076693667, - 0.006646841630),
    to_complex(- 0.013118414541, - 0.016413521278),
    to_complex(0.011334921437, - 0.000762369892),
    to_complex(0.006609443093, - 0.000419978586),
    to_complex(- 0.016392164168, - 0.020482027060),
    to_complex(0.079383226444, - 0.006725381148),
    to_complex(0.010007860539, - 0.003600022449),
    to_complex(- 0.082682399961, - 0.010900892666),
    to_complex(- 0.088458483369, - 0.011011451795),
    to_complex(0.016675767511, 0.063888125821),
    to_complex(0.000036374311, 0.028849766621),
    to_complex(0.018423165229, 0.007041295137),
    to_complex(0.020620057746, - 0.002701188546),
    to_complex(- 0.000215341506, - 0.030332046417),
    to_complex(0.032985823384, 0.019478447077),
    to_complex(- 0.018236706249, 0.044531009600),
    to_complex(0.046447866035, 0.025558954703),
    to_complex(0.021423875065, 0.077268929613),
    to_complex(0.063275623068, - 0.025830165752),
    to_complex(- 0.060530938589, - 0.066764397687),
    to_complex(0.103002651867, 0.038400767017),
    to_complex(0.014354195116, 0.083525752387),
    to_complex(- 0.022397016649, - 0.054292590786),
    to_complex(- 0.057900280945, - 0.129616093965),
    to_complex(- 0.039677687738, 0.049124724091),
    to_complex(- 0.001102295331, - 0.010727735201),
    to_complex(0.016935883028, 0.039871122307),
    to_complex(- 0.034332743850, 0.056996841989),
    to_complex(0.026637994948, 0.113442218433),
    to_complex(0.000734073926, 0.062729324104),
    to_complex(- 0.050653844489, 0.003910323478),
    to_complex(0.008691225801, 0.084426791615),
    to_complex(0.000612587631, - 0.002638110709),
    to_complex(0.015898052919, 0.039999066210),
    to_complex(0.048774305666, 0.019212382187),
    to_complex(0.071120771497, 0.017701851308),
    to_complex(0.082699026350, - 0.051118933877),
    to_complex(0.008512271530, - 0.051261741526),
    to_complex(- 0.061952733155, - 0.043820261007),
    to_complex(- 0.004449946878, 0.018600782532),
    to_complex(0.007349366365, 0.024865783526),
    to_complex(- 0.034405843202, 0.065531406366),
    to_complex(0.012924053117, 0.032784143524),
    to_complex(- 0.030686976264, - 0.005306035425),
    to_complex(- 0.034757430173, - 0.020383319961),
    to_complex(- 0.026895769223, - 0.013181349576),
    to_complex(0.094167600757, - 0.024741489636),
    to_complex(- 0.033951535470, 0.036977203566),
    to_complex(0.096488803983, 0.053746324123),
    to_complex(0.090556600363, - 0.021224217891),
    to_complex(0.019266854497, 0.018853380349),
    to_complex(0.060859515477, 0.033578979410),
    to_complex(- 0.021683278002, - 0.016722913910),
    to_complex(0.030270442666, - 0.120648781958),
    to_complex(0.034752457452, 0.032959303731),
    to_complex(- 0.024845901999, 0.071886208070),
    to_complex(- 0.047537345663, 0.053720869121),
    to_complex(- 0.045320384609, - 0.026559460967),
    to_complex(0.012603749187, 0.017107681541),
    to_complex(0.011211739557, - 0.044619960413),
    to_complex(0.043652152429, - 0.059172350354),
    to_complex(0.032733339395, - 0.018350916493),
    to_complex(0.083107483367, - 0.080044065416),
    to_complex(- 0.045607352973, 0.137898775589),
    to_complex(- 0.036518829038, 0.003028158051),
    to_complex(0.069445370405, - 0.054793157762),
    to_complex(0.022767172850, 0.080825449201),
    to_complex(0.001722347793, - 0.019010953469),
    to_complex(- 0.083310796657, - 0.044279882244),
    to_complex(0.099867503654, 0.058798059604),
    to_complex(0.027626670474, 0.021647778457),
    to_complex(0.050201913560, - 0.086054355247),
    to_complex(0.012005668902, 0.092462414438),
    to_complex(- 0.005586255035, - 0.029758962373),
    to_complex(- 0.000182239185, 0.009403743822),
    to_complex(- 0.061401572654, - 0.012807443943),
    to_complex(- 0.053339569330, - 0.008652440482),
    to_complex(0.029155656108, 0.051865218145),
    to_complex(- 0.020639707801, 0.045845872735),
    to_complex(0.083893418093, - 0.010501190332),
    to_complex(0.024632780871, 0.044161127942),
    to_complex(0.018436129763, 0.000704196592),
    to_complex(- 0.065598426004, 0.082739013885),
    to_complex(- 0.058725913897, - 0.096348738050),
    to_complex(- 0.000009930732, 0.111289881664),
    to_complex(- 0.053140496905, - 0.008768563987),
    to_complex(0.001560881716, - 0.055834666224),
    to_complex(0.001283937258, - 0.005889982909),
    to_complex(0.045259439376, - 0.065536563906),
    to_complex(0.002451210332, 0.035761477231),
    to_complex(- 0.042245257818, 0.002247978321),
    to_complex(- 0.032552872216, - 0.028068787522),
    to_complex(- 0.031819119684, - 0.086438178864),
    to_complex(- 0.007655114179, - 0.001856382892),
    to_complex(- 0.019422301116, - 0.100177732169),
    to_complex(0.017818752890, 0.015135475392),
    to_complex(0.025533064639, - 0.011307312964),
    to_complex(0.074675892098, - 0.059047770709),
    to_complex(0.015540511682, - 0.062221632481),
    to_complex(0.076372383861, - 0.034747237745),
    to_complex(- 0.028016358557, - 0.011672618920),
    to_complex(- 0.088444830971, - 0.009405296470),
    to_complex(0.012008407725, 0.004771150347),
    to_complex(0.045248326371, - 0.035044854165),
    to_complex(0.016989347252, - 0.007468152223),
    to_complex(0.028934464266, - 0.002391404184),
    to_complex(0.004809556586, - 0.031015116238),
    to_complex(- 0.024238375910, - 0.022229815312),
    to_complex(0.069212536383, - 0.085787334741),
    to_complex(0.037722852906, 0.029524049547),
    to_complex(0.157487546715, - 0.066240947701),
    to_complex(0.118844280294, - 0.062591248574),
    to_complex(- 0.023117034979, 0.053279790941),
    to_complex(- 0.059946741049, 0.006849783915),
    to_complex(- 0.000139550163, 0.035892693324),
    to_complex(- 0.043265070634, - 0.003800868047),
    to_complex(0.031800843331, - 0.053594918572),
    to_complex(0.025663674168, 0.019755637567),
    to_complex(- 0.018591833796, 0.035036314511),
    to_complex(0.059349186039, 0.063582149637),
    to_complex(0.054633630350, 0.102881018673),
    to_complex(- 0.044812164974, 0.037056906617),
    to_complex(0.078633737213, - 0.021764774796),
    to_complex(- 0.011218389041, 0.013510835918),
    to_complex(- 0.032126425385, - 0.029463964457),
    to_complex(- 0.069863173719, - 0.031184667409),
    to_complex(0.025613111539, - 0.010315012240),
    to_complex(0.057428584782, 0.068626022344),
    to_complex(- 0.041024181959, - 0.073304421272),
    to_complex(0.000213038732, - 0.010569088055),
    to_complex(0.018381500668, 0.043973803633),
    to_complex(0.097881200845, 0.011695094451),
    to_complex(- 0.048690680334, 0.028643069125),
    to_complex(- 0.037844590063, - 0.004242733484),
    to_complex(0.043931018499, - 0.030829287700),
    to_complex(0.012689526298, - 0.080093092855),
    to_complex(0.030065478730, - 0.005472140999),
    to_complex(- 0.036254332032, 0.150582598016),
    to_complex(- 0.010109024417, 0.059215550852),
    to_complex(- 0.047287815568, - 0.010744773116),
    to_complex(- 0.042981168370, 0.024439753120),
    to_complex(- 0.058048259373, 0.064685757190),
    to_complex(- 0.016175389924, 0.010378012531),
    to_complex(- 0.035650531562, 0.019666421696),
    to_complex(0.006105536778, - 0.063107981156),
    to_complex(- 0.104749432353, 0.068571151861),
    to_complex(- 0.039172325826, 0.002469533503),
    to_complex(- 0.041964983546, 0.048135156600),
    to_complex(- 0.010910246333, - 0.003931225343),
    to_complex(- 0.076020538639, - 0.033809193812),
    to_complex(- 0.005589291237, 0.101880043550),
    to_complex(0.008718486452, 0.033522174190),
    to_complex(0.087527162602, - 0.016311719380),
    to_complex(0.034939993226, 0.023314167717),
    to_complex(0.046498549360, - 0.007557256839),
    to_complex(0.040582800635, 0.005962319213),
    to_complex(- 0.015311702205, - 0.095376204475),
    to_complex(0.039142334444, 0.093518159435),
    to_complex(0.084653064739, 0.011900919266),
    to_complex(- 0.087366792246, - 0.011327777274),
    to_complex(0.003585835908, 0.026899677355),
    to_complex(- 0.033336006759, - 0.053488216865),
    to_complex(- 0.034344465195, 0.093574198807),
    to_complex(- 0.034556355364, 0.006865228050),
    to_complex(- 0.031740589896, 0.005949095074),
    to_complex(- 0.042536327163, - 0.042004556864),
    to_complex(- 0.006083670127, - 0.046151104784),
    to_complex(0.015993198488, 0.014349912009),
    to_complex(0.056711833461, - 0.008134046955),
    to_complex(0.036095755779, - 0.008297373653),
    to_complex(- 0.070566570297, - 0.013612973845),
    to_complex(- 0.041712828336, 0.044523574960),
    to_complex(0.054936682576, - 0.010392156504),
    to_complex(- 0.011271724619, 0.082782198532),
    to_complex(- 0.073324744949, 0.061462076215),
    to_complex(- 0.025588206764, - 0.013442203296),
    to_complex(0.000444371895, 0.064693652917),
    to_complex(- 0.064948198257, 0.029750715696),
    to_complex(0.054374886302, - 0.025527679057),
    to_complex(0.117355059675, - 0.048176367391),
    to_complex(- 0.004262159094, - 0.058156197372),
    to_complex(- 0.042252712953, - 0.020772986252),
    to_complex(0.052105600240, - 0.014474609251),
    to_complex(- 0.065585450820, - 0.006441152486),
    to_complex(- 0.089556506290, 0.036912635098),
    to_complex(0.019686412427, - 0.013340962240),
    to_complex(- 0.045893190675, - 0.023276498419),
    to_complex(0.017558621267, - 0.060752146768),
    to_complex(0.002940744699, 0.002567831274),
    to_complex(0.018173884007, 0.023368312249),
    to_complex(- 0.054875143838, 0.025004162570),
    to_complex(- 0.014087742971, 0.044740409114),
    to_complex(0.035887215602, 0.007905363739),
    to_complex(- 0.014413294988, 0.064730070955),
    to_complex(- 0.003052875676, 0.099128242713),
    to_complex(- 0.082714833286, - 0.094652550491),
    to_complex(0.053674332414, 0.064137282971),
    to_complex(0.034734003764, - 0.016225817075),
    to_complex(- 0.026872444646, - 0.055271282064),
    to_complex(0.027318670138, - 0.059066052548),
    to_complex(0.009715409320, 0.030866275522),
    to_complex(- 0.049013826033, 0.011636884523),
    to_complex(- 0.068369406042, - 0.038992922730),
    to_complex(0.043784599591, 0.017961436521),
    to_complex(- 0.080442613782, 0.017320570463),
    to_complex(- 0.012460807348, 0.063269089379),
    to_complex(0.095430067726, 0.096040316941),
    to_complex(0.058272099442, 0.047734973108),
    to_complex(- 0.057246447689, - 0.017470557604),
    to_complex(- 0.002635412386, 0.034023850119),
    to_complex(0.040168290250, 0.026693656665),
    to_complex(0.127290747991, - 0.019689552456),
    to_complex(- 0.017005877514, - 0.003012506793),
    to_complex(- 0.070067835935, - 0.016964486248),
    to_complex(0.023373891227, 0.082887697724),
    to_complex(0.037526417655, - 0.018819063780),
    to_complex(0.011179564537, 0.001695470785),
    to_complex(0.032366267204, - 0.079067732999),
    to_complex(- 0.107260896858, - 0.028523084834),
    to_complex(0.030693442276, - 0.060753940429),
    to_complex(- 0.016068638767, - 0.017995413808),
    to_complex(0.008790839545, - 0.099490937274),
    to_complex(- 0.057393492673, - 0.015800113714),
    to_complex(0.014839481961, - 0.018452237701),
    to_complex(0.124258518792, - 0.064811568171),
    to_complex(- 0.024508442648, - 0.065202456305),
    to_complex(- 0.041192418953, 0.006540452644),
    to_complex(0.003775274680, 0.039772476168),
    to_complex(- 0.127813117082, - 0.022529086205),
    to_complex(0.011093604751, 0.005510893265),
    to_complex(- 0.064799604370, - 0.072838254494),
    to_complex(- 0.061335612863, - 0.015338911038),
    to_complex(0.000700373816, 0.015555567322),
    to_complex(0.046328646002, 0.029679802029),
    to_complex(0.073283831110, - 0.056531909538),
    to_complex(- 0.039295378169, 0.009561765859),
    to_complex(0.058607522960, - 0.020454292234),
    to_complex(0.043176068873, - 0.097745936845),
    to_complex(0.027410111904, - 0.022901785461),
    to_complex(- 0.050624956278, - 0.005470003482),
    to_complex(- 0.085056162099, 0.046986226834),
    to_complex(- 0.026295056500, 0.020886120758),
    to_complex(0.068227219035, 0.046988682955),
    to_complex(0.039559723436, - 0.023076353306),
    to_complex(0.024521174130, - 0.068245273230),
    to_complex(- 0.033452288242, - 0.033294503408),
    to_complex(0.085205156248, 0.017065071121),
    to_complex(- 0.014689238363, 0.034415456859),
    to_complex(0.010117101951, 0.004684447377),
    to_complex(0.025196704313, - 0.033712851193),
    to_complex(- 0.009478758482, 0.003993353853),
    to_complex(- 0.047982603977, 0.087210214675),
    to_complex(- 0.047611723807, - 0.016086658258),
    to_complex(- 0.059040348920, 0.017393852270),
    to_complex(- 0.060211191748, - 0.041742575421),
    to_complex(0.018535971361, - 0.005718885441),
    to_complex(- 0.040487899459, - 0.047311005694),
    to_complex(0.002456149958, 0.052719380946),
    to_complex(0.036351263033, 0.039140744994),
    to_complex(- 0.058656651729, 0.001039467198),
    to_complex(- 0.059900805459, 0.022679600056),
    to_complex(- 0.001704654174, 0.018437717147),
    to_complex(0.028727796180, 0.083423582693),
    to_complex(- 0.084338532405, 0.072083207875),
    to_complex(- 0.008786815540, - 0.007543510775),
    to_complex(0.004575786896, - 0.072670901641),
    to_complex(0.006469711556, - 0.047868238122),
    to_complex(0.028416931955, 0.095875034249),
    to_complex(- 0.097766386455, - 0.156380938193),
    to_complex(0.021814270117, 0.035709621966),
    to_complex(- 0.020697284325, 0.120448946973),
    to_complex(- 0.029175899506, - 0.034036807077),
    to_complex(0.052430672852, - 0.001446228779),
    to_complex(- 0.030357849134, 0.001656527387),
    to_complex(- 0.025394555425, - 0.011072477755),
    to_complex(0.013022861879, - 0.034906195588),
    to_complex(0.074519856818, 0.031877632206),
    to_complex(- 0.105438269973, 0.006433141240),
    to_complex(0.053072392772, - 0.010300222945),
    to_complex(- 0.070589864334, - 0.028392416666),
    to_complex(0.027378868056, 0.042264555167),
    to_complex(0.078738513562, - 0.071353376456),
    to_complex(0.057707375747, 0.003199629344),
    to_complex(0.072182921334, 0.031051097051),
    to_complex(- 0.034577966405, - 0.015001055286),
    to_complex(- 0.061832287190, 0.014613715133),
    to_complex(- 0.011814783926, - 0.050185714875),
    to_complex(- 0.070539453440, 0.083118958125),
    to_complex(0.057265823538, 0.028804110923),
    to_complex(- 0.043410473537, 0.027530572337),
    to_complex(0.042793875606, - 0.064876223880),
    to_complex(0.013162184537, 0.010614197365),
    to_complex(0.046936440120, 0.037571449199),
    to_complex(0.018515282655, - 0.084916531356),
    to_complex(- 0.009100786419, - 0.085119464790),
    to_complex(0.019889569006, - 0.021877209891),
    to_complex(- 0.031248570981, - 0.031543857797),
    to_complex(0.122893398776, 0.019954740641),
    to_complex(0.061318390798, 0.051174566893),
    to_complex(- 0.079080284354, 0.012921383978),
    to_complex(- 0.199251012075, - 0.051539615747),
    to_complex(0.041917898440, - 0.057548142233),
    to_complex(0.003338093970, 0.014072815880),
    to_complex(- 0.049286544921, - 0.034331268199),
    to_complex(- 0.022900224780, - 0.025389071376),
    to_complex(0.046044782562, 0.027152106448),
    to_complex(0.056973819827, - 0.067137580923),
    to_complex(0.005543124876, 0.041912841953),
    to_complex(- 0.072861093600, - 0.002512409654),
    to_complex(0.082338390751, 0.029980857799),
    to_complex(0.058323394075, - 0.020786867070),
    to_complex(- 0.050913812004, 0.055973734863),
    to_complex(- 0.067641226059, 0.026964337761),
    to_complex(- 0.002359424747, - 0.067827237835),
    to_complex(- 0.037389646327, - 0.026890781353),
    to_complex(- 0.109340907521, 0.021692890182),
    to_complex(0.007434102849, - 0.064728801036),
    to_complex(0.085329755074, - 0.072102805945),
    to_complex(0.025392617692, 0.031637836205),
    to_complex(0.004417591185, - 0.004054164803),
    to_complex(- 0.044211416228, - 0.018920879169),
    to_complex(- 0.048048929134, - 0.096586830997),
    to_complex(0.013910898217, 0.017774301955),
    to_complex(- 0.028618802296, 0.064196891430),
    to_complex(- 0.043266237299, 0.106487707480),
    to_complex(0.060767866413, 0.010116009281),
    to_complex(0.053676272635, 0.013603164501),
    to_complex(- 0.057322260965, - 0.059234341478),
    to_complex(0.030533220197, 0.071639772528),
    to_complex(0.028390615167, - 0.059518681379),
    to_complex(0.016887847944, - 0.080747548287),
    to_complex(0.020114421706, 0.045820888361),
    to_complex(- 0.037324091537, - 0.020927751918),
    to_complex(- 0.015962629490, 0.036331309601),
    to_complex(0.051663358461, 0.001962440197),
    to_complex(0.052196265883, - 0.018549303478),
    to_complex(0.042810070696, - 0.007392097739),
    to_complex(- 0.020375263717, 0.082404860759),
    to_complex(0.039097351231, - 0.026184365681),
    to_complex(- 0.002349194488, 0.020205863730),
    to_complex(- 0.085973526388, 0.054042862041),
    to_complex(- 0.024617946903, 0.022910693216),
    to_complex(- 0.000536126058, - 0.084069785812),
    to_complex(- 0.004004314682, 0.103951059225),
    to_complex(- 0.010747232794, - 0.081956006208),
    to_complex(0.010757078585, - 0.085363151282),
    to_complex(- 0.053115404741, 0.009622380263),
    to_complex(- 0.066493249336, 0.008786809901),
    to_complex(0.020909036281, 0.038371174920),
    to_complex(0.054672877930, 0.007770307919),
    to_complex(- 0.014933700788, - 0.049933595348),
    to_complex(0.047477120851, 0.030094236619),
    to_complex(- 0.079699434885, 0.083644752860),
    to_complex(0.142717329775, - 0.061564633162),
    to_complex(0.005354600473, 0.036177308147),
    to_complex(0.056815496599, - 0.009658548144),
    to_complex(0.050256699890, 0.033517798828),
    to_complex(- 0.043575742079, - 0.051386825533),
    to_complex(- 0.025373604772, 0.007733108674),
    to_complex(0.026667793180, - 0.041669878233),
    to_complex(0.013530707019, 0.007472720229),
    to_complex(- 0.008460512348, - 0.059503226059),
    to_complex(0.023811812169, - 0.071946737576),
    to_complex(0.050706892360, - 0.047585317899),
    to_complex(0.006698542688, - 0.084384750039),
    to_complex(0.033456826051, - 0.010139577192),
    to_complex(0.040584794729, - 0.025662869228),
    to_complex(0.009072570592, 0.033416780851),
    to_complex(- 0.093377416404, - 0.002614579166),
    to_complex(- 0.033706949066, - 0.033138226497),
    to_complex(- 0.024245084285, 0.026034113293),
    to_complex(0.015440111890, 0.063382986277),
    to_complex(- 0.052737332390, - 0.160082011744),
    to_complex(0.123942968927, 0.012015604732),
    to_complex(0.041543226871, 0.017030255611),
    to_complex(- 0.014434840602, - 0.045976523797),
    to_complex(0.014655931546, 0.000333626344),
    to_complex(- 0.055079668215, 0.004061737072),
    to_complex(0.043875284087, - 0.067691436247),
    to_complex(0.079373239861, - 0.088948313635),
    to_complex(- 0.031731362471, 0.021239613240),
    to_complex(- 0.020850857206, 0.015004298003),
    to_complex(0.038299319274, 0.035249787192),
    to_complex(0.112228806761, 0.029947801219),
    to_complex(0.013706063617, 0.027344895795),
    to_complex(0.041957499476, - 0.010862535372),
    to_complex(- 0.068184301884, 0.074203458021),
    to_complex(- 0.048315749132, 0.018728904080),
    to_complex(- 0.022704147366, - 0.073484546079),
    to_complex(0.006926829731, - 0.036390485790),
    to_complex(- 0.025077991064, 0.081992607068),
    to_complex(0.018974978108, 0.054318144781),
    to_complex(0.001056478747, 0.014182360632),
    to_complex(0.046006979074, - 0.066290429833),
    to_complex(- 0.000043426526, 0.019632249214),
    to_complex(- 0.046848498433, - 0.012621373025),
    to_complex(0.004034284890, 0.010022385852),
    to_complex(- 0.058894251216, 0.012390728329),
    to_complex(- 0.046917073501, - 0.088308636848),
    to_complex(- 0.016508147056, 0.002457591251),
    to_complex(- 0.018818866105, - 0.042779702005),
    to_complex(0.058067487154, 0.017190002489),
    to_complex(- 0.047883419853, - 0.051687214522),
    to_complex(- 0.020252589887, - 0.015557542400),
    to_complex(- 0.052377412058, - 0.025378605838),
    to_complex(- 0.100541216675, 0.133907914960),
    to_complex(- 0.051846423473, - 0.011141584790),
    to_complex(- 0.095504417956, 0.086516011009),
    to_complex(0.049531876683, - 0.045247897683),
    to_complex(0.051477955532, 0.080880411375),
    to_complex(0.037643107603, - 0.039985208680),
    to_complex(0.019027570855, - 0.099743049475),
    to_complex(- 0.032468252651, 0.007574273285),
    to_complex(- 0.075702695219, 0.038535919031),
    to_complex(- 0.090339341444, 0.039615424118),
    to_complex(- 0.051081425014, 0.048445238190),
    to_complex(0.007992929276, 0.018433665211),
    to_complex(0.014029930307, 0.002938679038),
    to_complex(0.069547729966, - 0.071949617751),
    to_complex(- 0.063017614991, - 0.022669916979),
    to_complex(0.000817181094, - 0.067287914199),
    to_complex(0.020385600417, 0.062256091161),
    to_complex(0.066917078363, 0.012347076617),
    to_complex(- 0.083112825668, - 0.038305054147),
    to_complex(- 0.006956041053, - 0.004641267003),
    to_complex(0.047736611147, 0.096582113905),
    to_complex(0.026069253728, 0.012455746506),
    to_complex(- 0.041257833168, 0.002019150236),
    to_complex(0.022032840361, 0.047662666173),
    to_complex(0.007562896646, - 0.097667143103),
    to_complex(- 0.025402012929, 0.018617027701),
    to_complex(0.036880709730, - 0.009612289745),
    to_complex(- 0.012726896802, 0.030693076600),
    to_complex(0.089667541108, - 0.014273106537),
    to_complex(0.034055454096, - 0.012724509042),
    to_complex(- 0.080162050700, 0.069534950889),
    to_complex(- 0.069543994699, 0.004168591600),
    to_complex(0.040477320552, 0.022139282577),
    to_complex(0.052033213583, - 0.070088240450),
    to_complex(- 0.047545581228, 0.007008703862),
    to_complex(- 0.015774581627, - 0.065494577664),
    to_complex(0.016901632439, - 0.057824790988),
    to_complex(- 0.054234621557, - 0.076556239018),
    to_complex(- 0.053800708793, - 0.063581214027),
    to_complex(0.024688264008, 0.022209193867),
    to_complex(0.013276874429, - 0.097258275183),
    to_complex(- 0.031415933193, - 0.021935943450),
    to_complex(- 0.045214279159, 0.039216112171),
    to_complex(0.091327555991, 0.040439653587),
    to_complex(- 0.008024007099, - 0.000954114002),
    to_complex(0.081902677377, 0.004242049439),
    to_complex(0.027322180892, 0.122579128793),
    to_complex(- 0.052874078633, - 0.067296246592),
    to_complex(- 0.049732049753, 0.037227685604));

end package;
