library IEEE;
  use work.complex_pkg.all;

package twiddle_values is

  constant TWIDDLE_VALUES_2048 : complex_array(0 to 1023) := (
    to_complex(1.000000000000, 0.000000000000),
    to_complex(1.000000000000, - 0.003173828125),
    to_complex(1.000000000000, - 0.006103515625),
    to_complex(1.000000000000, - 0.009277343750),
    to_complex(1.000000000000, - 0.012207031250),
    to_complex(1.000000000000, - 0.015380859375),
    to_complex(0.999755859375, - 0.018310546875),
    to_complex(0.999755859375, - 0.021484375000),
    to_complex(0.999755859375, - 0.024658203125),
    to_complex(0.999511718750, - 0.027587890625),
    to_complex(0.999511718750, - 0.030761718750),
    to_complex(0.999511718750, - 0.033691406250),
    to_complex(0.999267578125, - 0.036865234375),
    to_complex(0.999267578125, - 0.039794921875),
    to_complex(0.999023437500, - 0.042968750000),
    to_complex(0.999023437500, - 0.045898437500),
    to_complex(0.998779296875, - 0.049072265625),
    to_complex(0.998535156250, - 0.052246093750),
    to_complex(0.998535156250, - 0.055175781250),
    to_complex(0.998291015625, - 0.058349609375),
    to_complex(0.998046875000, - 0.061279296875),
    to_complex(0.998046875000, - 0.064453125000),
    to_complex(0.997802734375, - 0.067382812500),
    to_complex(0.997558593750, - 0.070556640625),
    to_complex(0.997314453125, - 0.073486328125),
    to_complex(0.997070312500, - 0.076660156250),
    to_complex(0.996826171875, - 0.079589843750),
    to_complex(0.996582031250, - 0.082763671875),
    to_complex(0.996337890625, - 0.085693359375),
    to_complex(0.996093750000, - 0.088867187500),
    to_complex(0.995849609375, - 0.091796875000),
    to_complex(0.995361328125, - 0.094970703125),
    to_complex(0.995117187500, - 0.097900390625),
    to_complex(0.994873046875, - 0.101074218750),
    to_complex(0.994628906250, - 0.104003906250),
    to_complex(0.994140625000, - 0.107177734375),
    to_complex(0.993896484375, - 0.110107421875),
    to_complex(0.993652343750, - 0.113281250000),
    to_complex(0.993164062500, - 0.116210937500),
    to_complex(0.992919921875, - 0.119384765625),
    to_complex(0.992431640625, - 0.122314453125),
    to_complex(0.992187500000, - 0.125488281250),
    to_complex(0.991699218750, - 0.128417968750),
    to_complex(0.991210937500, - 0.131591796875),
    to_complex(0.990966796875, - 0.134521484375),
    to_complex(0.990478515625, - 0.137695312500),
    to_complex(0.989990234375, - 0.140625000000),
    to_complex(0.989501953125, - 0.143798828125),
    to_complex(0.989257812500, - 0.146728515625),
    to_complex(0.988769531250, - 0.149658203125),
    to_complex(0.988281250000, - 0.152832031250),
    to_complex(0.987792968750, - 0.155761718750),
    to_complex(0.987304687500, - 0.158935546875),
    to_complex(0.986816406250, - 0.161865234375),
    to_complex(0.986328125000, - 0.164794921875),
    to_complex(0.985839843750, - 0.167968750000),
    to_complex(0.985351562500, - 0.170898437500),
    to_complex(0.984863281250, - 0.174072265625),
    to_complex(0.984130859375, - 0.177001953125),
    to_complex(0.983642578125, - 0.179931640625),
    to_complex(0.983154296875, - 0.183105468750),
    to_complex(0.982421875000, - 0.186035156250),
    to_complex(0.981933593750, - 0.188964843750),
    to_complex(0.981445312500, - 0.192138671875),
    to_complex(0.980712890625, - 0.195068359375),
    to_complex(0.980224609375, - 0.197998046875),
    to_complex(0.979492187500, - 0.201171875000),
    to_complex(0.979003906250, - 0.204101562500),
    to_complex(0.978271484375, - 0.207031250000),
    to_complex(0.977783203125, - 0.210205078125),
    to_complex(0.977050781250, - 0.213134765625),
    to_complex(0.976318359375, - 0.216064453125),
    to_complex(0.975585937500, - 0.218994140625),
    to_complex(0.975097656250, - 0.222167968750),
    to_complex(0.974365234375, - 0.225097656250),
    to_complex(0.973632812500, - 0.228027343750),
    to_complex(0.972900390625, - 0.230957031250),
    to_complex(0.972167968750, - 0.234130859375),
    to_complex(0.971435546875, - 0.237060546875),
    to_complex(0.970703125000, - 0.239990234375),
    to_complex(0.969970703125, - 0.242919921875),
    to_complex(0.969238281250, - 0.245849609375),
    to_complex(0.968505859375, - 0.249023437500),
    to_complex(0.967773437500, - 0.251953125000),
    to_complex(0.967041015625, - 0.254882812500),
    to_complex(0.966308593750, - 0.257812500000),
    to_complex(0.965332031250, - 0.260742187500),
    to_complex(0.964599609375, - 0.263671875000),
    to_complex(0.963867187500, - 0.266601562500),
    to_complex(0.962890625000, - 0.269775390625),
    to_complex(0.962158203125, - 0.272705078125),
    to_complex(0.961181640625, - 0.275634765625),
    to_complex(0.960449218750, - 0.278564453125),
    to_complex(0.959472656250, - 0.281494140625),
    to_complex(0.958740234375, - 0.284423828125),
    to_complex(0.957763671875, - 0.287353515625),
    to_complex(0.957031250000, - 0.290283203125),
    to_complex(0.956054687500, - 0.293212890625),
    to_complex(0.955078125000, - 0.296142578125),
    to_complex(0.954345703125, - 0.299072265625),
    to_complex(0.953369140625, - 0.302001953125),
    to_complex(0.952392578125, - 0.304931640625),
    to_complex(0.951416015625, - 0.307861328125),
    to_complex(0.950439453125, - 0.310791015625),
    to_complex(0.949462890625, - 0.313720703125),
    to_complex(0.948486328125, - 0.316650390625),
    to_complex(0.947509765625, - 0.319580078125),
    to_complex(0.946533203125, - 0.322509765625),
    to_complex(0.945556640625, - 0.325195312500),
    to_complex(0.944580078125, - 0.328125000000),
    to_complex(0.943603515625, - 0.331054687500),
    to_complex(0.942626953125, - 0.333984375000),
    to_complex(0.941650390625, - 0.336914062500),
    to_complex(0.940429687500, - 0.339843750000),
    to_complex(0.939453125000, - 0.342773437500),
    to_complex(0.938476562500, - 0.345458984375),
    to_complex(0.937255859375, - 0.348388671875),
    to_complex(0.936279296875, - 0.351318359375),
    to_complex(0.935302734375, - 0.354248046875),
    to_complex(0.934082031250, - 0.356933593750),
    to_complex(0.933105468750, - 0.359863281250),
    to_complex(0.931884765625, - 0.362792968750),
    to_complex(0.930664062500, - 0.365722656250),
    to_complex(0.929687500000, - 0.368408203125),
    to_complex(0.928466796875, - 0.371337890625),
    to_complex(0.927246093750, - 0.374267578125),
    to_complex(0.926269531250, - 0.376953125000),
    to_complex(0.925048828125, - 0.379882812500),
    to_complex(0.923828125000, - 0.382568359375),
    to_complex(0.922607421875, - 0.385498046875),
    to_complex(0.921630859375, - 0.388427734375),
    to_complex(0.920410156250, - 0.391113281250),
    to_complex(0.919189453125, - 0.394042968750),
    to_complex(0.917968750000, - 0.396728515625),
    to_complex(0.916748046875, - 0.399658203125),
    to_complex(0.915527343750, - 0.402343750000),
    to_complex(0.914306640625, - 0.405273437500),
    to_complex(0.912841796875, - 0.407958984375),
    to_complex(0.911621093750, - 0.410888671875),
    to_complex(0.910400390625, - 0.413574218750),
    to_complex(0.909179687500, - 0.416503906250),
    to_complex(0.907958984375, - 0.419189453125),
    to_complex(0.906494140625, - 0.422119140625),
    to_complex(0.905273437500, - 0.424804687500),
    to_complex(0.904052734375, - 0.427490234375),
    to_complex(0.902587890625, - 0.430419921875),
    to_complex(0.901367187500, - 0.433105468750),
    to_complex(0.899902343750, - 0.435791015625),
    to_complex(0.898681640625, - 0.438720703125),
    to_complex(0.897216796875, - 0.441406250000),
    to_complex(0.895996093750, - 0.444091796875),
    to_complex(0.894531250000, - 0.446777343750),
    to_complex(0.893310546875, - 0.449707031250),
    to_complex(0.891845703125, - 0.452392578125),
    to_complex(0.890380859375, - 0.455078125000),
    to_complex(0.889160156250, - 0.457763671875),
    to_complex(0.887695312500, - 0.460449218750),
    to_complex(0.886230468750, - 0.463378906250),
    to_complex(0.884765625000, - 0.466064453125),
    to_complex(0.883300781250, - 0.468750000000),
    to_complex(0.881835937500, - 0.471435546875),
    to_complex(0.880371093750, - 0.474121093750),
    to_complex(0.878906250000, - 0.476806640625),
    to_complex(0.877441406250, - 0.479492187500),
    to_complex(0.875976562500, - 0.482177734375),
    to_complex(0.874511718750, - 0.484863281250),
    to_complex(0.873046875000, - 0.487548828125),
    to_complex(0.871582031250, - 0.490234375000),
    to_complex(0.870117187500, - 0.492919921875),
    to_complex(0.868652343750, - 0.495605468750),
    to_complex(0.866943359375, - 0.498291015625),
    to_complex(0.865478515625, - 0.500976562500),
    to_complex(0.864013671875, - 0.503417968750),
    to_complex(0.862304687500, - 0.506103515625),
    to_complex(0.860839843750, - 0.508789062500),
    to_complex(0.859375000000, - 0.511474609375),
    to_complex(0.857666015625, - 0.514160156250),
    to_complex(0.856201171875, - 0.516845703125),
    to_complex(0.854492187500, - 0.519287109375),
    to_complex(0.853027343750, - 0.521972656250),
    to_complex(0.851318359375, - 0.524658203125),
    to_complex(0.849853515625, - 0.527099609375),
    to_complex(0.848144531250, - 0.529785156250),
    to_complex(0.846435546875, - 0.532470703125),
    to_complex(0.844970703125, - 0.534912109375),
    to_complex(0.843261718750, - 0.537597656250),
    to_complex(0.841552734375, - 0.540283203125),
    to_complex(0.839843750000, - 0.542724609375),
    to_complex(0.838134765625, - 0.545410156250),
    to_complex(0.836425781250, - 0.547851562500),
    to_complex(0.834960937500, - 0.550537109375),
    to_complex(0.833251953125, - 0.552978515625),
    to_complex(0.831542968750, - 0.555664062500),
    to_complex(0.829833984375, - 0.558105468750),
    to_complex(0.828125000000, - 0.560546875000),
    to_complex(0.826416015625, - 0.563232421875),
    to_complex(0.824707031250, - 0.565673828125),
    to_complex(0.822753906250, - 0.568359375000),
    to_complex(0.821044921875, - 0.570800781250),
    to_complex(0.819335937500, - 0.573242187500),
    to_complex(0.817626953125, - 0.575927734375),
    to_complex(0.815917968750, - 0.578369140625),
    to_complex(0.813964843750, - 0.580810546875),
    to_complex(0.812255859375, - 0.583251953125),
    to_complex(0.810546875000, - 0.585693359375),
    to_complex(0.808593750000, - 0.588378906250),
    to_complex(0.806884765625, - 0.590820312500),
    to_complex(0.804931640625, - 0.593261718750),
    to_complex(0.803222656250, - 0.595703125000),
    to_complex(0.801269531250, - 0.598144531250),
    to_complex(0.799560546875, - 0.600585937500),
    to_complex(0.797607421875, - 0.603027343750),
    to_complex(0.795898437500, - 0.605468750000),
    to_complex(0.793945312500, - 0.607910156250),
    to_complex(0.791992187500, - 0.610351562500),
    to_complex(0.790283203125, - 0.612792968750),
    to_complex(0.788330078125, - 0.615234375000),
    to_complex(0.786376953125, - 0.617675781250),
    to_complex(0.784667968750, - 0.620117187500),
    to_complex(0.782714843750, - 0.622558593750),
    to_complex(0.780761718750, - 0.624755859375),
    to_complex(0.778808593750, - 0.627197265625),
    to_complex(0.776855468750, - 0.629638671875),
    to_complex(0.774902343750, - 0.632080078125),
    to_complex(0.772949218750, - 0.634277343750),
    to_complex(0.770996093750, - 0.636718750000),
    to_complex(0.769042968750, - 0.639160156250),
    to_complex(0.767089843750, - 0.641601562500),
    to_complex(0.765136718750, - 0.643798828125),
    to_complex(0.763183593750, - 0.646240234375),
    to_complex(0.761230468750, - 0.648437500000),
    to_complex(0.759277343750, - 0.650878906250),
    to_complex(0.757324218750, - 0.653076171875),
    to_complex(0.755126953125, - 0.655517578125),
    to_complex(0.753173828125, - 0.657714843750),
    to_complex(0.751220703125, - 0.660156250000),
    to_complex(0.749023437500, - 0.662353515625),
    to_complex(0.747070312500, - 0.664794921875),
    to_complex(0.745117187500, - 0.666992187500),
    to_complex(0.742919921875, - 0.669189453125),
    to_complex(0.740966796875, - 0.671630859375),
    to_complex(0.738769531250, - 0.673828125000),
    to_complex(0.736816406250, - 0.676025390625),
    to_complex(0.734619140625, - 0.678466796875),
    to_complex(0.732666015625, - 0.680664062500),
    to_complex(0.730468750000, - 0.682861328125),
    to_complex(0.728515625000, - 0.685058593750),
    to_complex(0.726318359375, - 0.687255859375),
    to_complex(0.724365234375, - 0.689453125000),
    to_complex(0.722167968750, - 0.691650390625),
    to_complex(0.719970703125, - 0.694091796875),
    to_complex(0.717773437500, - 0.696289062500),
    to_complex(0.715820312500, - 0.698486328125),
    to_complex(0.713623046875, - 0.700683593750),
    to_complex(0.711425781250, - 0.702636718750),
    to_complex(0.709228515625, - 0.704833984375),
    to_complex(0.707031250000, - 0.707031250000),
    to_complex(0.704833984375, - 0.709228515625),
    to_complex(0.702636718750, - 0.711425781250),
    to_complex(0.700683593750, - 0.713623046875),
    to_complex(0.698486328125, - 0.715820312500),
    to_complex(0.696289062500, - 0.717773437500),
    to_complex(0.694091796875, - 0.719970703125),
    to_complex(0.691650390625, - 0.722167968750),
    to_complex(0.689453125000, - 0.724365234375),
    to_complex(0.687255859375, - 0.726318359375),
    to_complex(0.685058593750, - 0.728515625000),
    to_complex(0.682861328125, - 0.730468750000),
    to_complex(0.680664062500, - 0.732666015625),
    to_complex(0.678466796875, - 0.734619140625),
    to_complex(0.676025390625, - 0.736816406250),
    to_complex(0.673828125000, - 0.738769531250),
    to_complex(0.671630859375, - 0.740966796875),
    to_complex(0.669189453125, - 0.742919921875),
    to_complex(0.666992187500, - 0.745117187500),
    to_complex(0.664794921875, - 0.747070312500),
    to_complex(0.662353515625, - 0.749023437500),
    to_complex(0.660156250000, - 0.751220703125),
    to_complex(0.657714843750, - 0.753173828125),
    to_complex(0.655517578125, - 0.755126953125),
    to_complex(0.653076171875, - 0.757324218750),
    to_complex(0.650878906250, - 0.759277343750),
    to_complex(0.648437500000, - 0.761230468750),
    to_complex(0.646240234375, - 0.763183593750),
    to_complex(0.643798828125, - 0.765136718750),
    to_complex(0.641601562500, - 0.767089843750),
    to_complex(0.639160156250, - 0.769042968750),
    to_complex(0.636718750000, - 0.770996093750),
    to_complex(0.634277343750, - 0.772949218750),
    to_complex(0.632080078125, - 0.774902343750),
    to_complex(0.629638671875, - 0.776855468750),
    to_complex(0.627197265625, - 0.778808593750),
    to_complex(0.624755859375, - 0.780761718750),
    to_complex(0.622558593750, - 0.782714843750),
    to_complex(0.620117187500, - 0.784667968750),
    to_complex(0.617675781250, - 0.786376953125),
    to_complex(0.615234375000, - 0.788330078125),
    to_complex(0.612792968750, - 0.790283203125),
    to_complex(0.610351562500, - 0.791992187500),
    to_complex(0.607910156250, - 0.793945312500),
    to_complex(0.605468750000, - 0.795898437500),
    to_complex(0.603027343750, - 0.797607421875),
    to_complex(0.600585937500, - 0.799560546875),
    to_complex(0.598144531250, - 0.801269531250),
    to_complex(0.595703125000, - 0.803222656250),
    to_complex(0.593261718750, - 0.804931640625),
    to_complex(0.590820312500, - 0.806884765625),
    to_complex(0.588378906250, - 0.808593750000),
    to_complex(0.585693359375, - 0.810546875000),
    to_complex(0.583251953125, - 0.812255859375),
    to_complex(0.580810546875, - 0.813964843750),
    to_complex(0.578369140625, - 0.815917968750),
    to_complex(0.575927734375, - 0.817626953125),
    to_complex(0.573242187500, - 0.819335937500),
    to_complex(0.570800781250, - 0.821044921875),
    to_complex(0.568359375000, - 0.822753906250),
    to_complex(0.565673828125, - 0.824707031250),
    to_complex(0.563232421875, - 0.826416015625),
    to_complex(0.560546875000, - 0.828125000000),
    to_complex(0.558105468750, - 0.829833984375),
    to_complex(0.555664062500, - 0.831542968750),
    to_complex(0.552978515625, - 0.833251953125),
    to_complex(0.550537109375, - 0.834960937500),
    to_complex(0.547851562500, - 0.836425781250),
    to_complex(0.545410156250, - 0.838134765625),
    to_complex(0.542724609375, - 0.839843750000),
    to_complex(0.540283203125, - 0.841552734375),
    to_complex(0.537597656250, - 0.843261718750),
    to_complex(0.534912109375, - 0.844970703125),
    to_complex(0.532470703125, - 0.846435546875),
    to_complex(0.529785156250, - 0.848144531250),
    to_complex(0.527099609375, - 0.849853515625),
    to_complex(0.524658203125, - 0.851318359375),
    to_complex(0.521972656250, - 0.853027343750),
    to_complex(0.519287109375, - 0.854492187500),
    to_complex(0.516845703125, - 0.856201171875),
    to_complex(0.514160156250, - 0.857666015625),
    to_complex(0.511474609375, - 0.859375000000),
    to_complex(0.508789062500, - 0.860839843750),
    to_complex(0.506103515625, - 0.862304687500),
    to_complex(0.503417968750, - 0.864013671875),
    to_complex(0.500976562500, - 0.865478515625),
    to_complex(0.498291015625, - 0.866943359375),
    to_complex(0.495605468750, - 0.868652343750),
    to_complex(0.492919921875, - 0.870117187500),
    to_complex(0.490234375000, - 0.871582031250),
    to_complex(0.487548828125, - 0.873046875000),
    to_complex(0.484863281250, - 0.874511718750),
    to_complex(0.482177734375, - 0.875976562500),
    to_complex(0.479492187500, - 0.877441406250),
    to_complex(0.476806640625, - 0.878906250000),
    to_complex(0.474121093750, - 0.880371093750),
    to_complex(0.471435546875, - 0.881835937500),
    to_complex(0.468750000000, - 0.883300781250),
    to_complex(0.466064453125, - 0.884765625000),
    to_complex(0.463378906250, - 0.886230468750),
    to_complex(0.460449218750, - 0.887695312500),
    to_complex(0.457763671875, - 0.889160156250),
    to_complex(0.455078125000, - 0.890380859375),
    to_complex(0.452392578125, - 0.891845703125),
    to_complex(0.449707031250, - 0.893310546875),
    to_complex(0.446777343750, - 0.894531250000),
    to_complex(0.444091796875, - 0.895996093750),
    to_complex(0.441406250000, - 0.897216796875),
    to_complex(0.438720703125, - 0.898681640625),
    to_complex(0.435791015625, - 0.899902343750),
    to_complex(0.433105468750, - 0.901367187500),
    to_complex(0.430419921875, - 0.902587890625),
    to_complex(0.427490234375, - 0.904052734375),
    to_complex(0.424804687500, - 0.905273437500),
    to_complex(0.422119140625, - 0.906494140625),
    to_complex(0.419189453125, - 0.907958984375),
    to_complex(0.416503906250, - 0.909179687500),
    to_complex(0.413574218750, - 0.910400390625),
    to_complex(0.410888671875, - 0.911621093750),
    to_complex(0.407958984375, - 0.912841796875),
    to_complex(0.405273437500, - 0.914306640625),
    to_complex(0.402343750000, - 0.915527343750),
    to_complex(0.399658203125, - 0.916748046875),
    to_complex(0.396728515625, - 0.917968750000),
    to_complex(0.394042968750, - 0.919189453125),
    to_complex(0.391113281250, - 0.920410156250),
    to_complex(0.388427734375, - 0.921630859375),
    to_complex(0.385498046875, - 0.922607421875),
    to_complex(0.382568359375, - 0.923828125000),
    to_complex(0.379882812500, - 0.925048828125),
    to_complex(0.376953125000, - 0.926269531250),
    to_complex(0.374267578125, - 0.927246093750),
    to_complex(0.371337890625, - 0.928466796875),
    to_complex(0.368408203125, - 0.929687500000),
    to_complex(0.365722656250, - 0.930664062500),
    to_complex(0.362792968750, - 0.931884765625),
    to_complex(0.359863281250, - 0.933105468750),
    to_complex(0.356933593750, - 0.934082031250),
    to_complex(0.354248046875, - 0.935302734375),
    to_complex(0.351318359375, - 0.936279296875),
    to_complex(0.348388671875, - 0.937255859375),
    to_complex(0.345458984375, - 0.938476562500),
    to_complex(0.342773437500, - 0.939453125000),
    to_complex(0.339843750000, - 0.940429687500),
    to_complex(0.336914062500, - 0.941650390625),
    to_complex(0.333984375000, - 0.942626953125),
    to_complex(0.331054687500, - 0.943603515625),
    to_complex(0.328125000000, - 0.944580078125),
    to_complex(0.325195312500, - 0.945556640625),
    to_complex(0.322509765625, - 0.946533203125),
    to_complex(0.319580078125, - 0.947509765625),
    to_complex(0.316650390625, - 0.948486328125),
    to_complex(0.313720703125, - 0.949462890625),
    to_complex(0.310791015625, - 0.950439453125),
    to_complex(0.307861328125, - 0.951416015625),
    to_complex(0.304931640625, - 0.952392578125),
    to_complex(0.302001953125, - 0.953369140625),
    to_complex(0.299072265625, - 0.954345703125),
    to_complex(0.296142578125, - 0.955078125000),
    to_complex(0.293212890625, - 0.956054687500),
    to_complex(0.290283203125, - 0.957031250000),
    to_complex(0.287353515625, - 0.957763671875),
    to_complex(0.284423828125, - 0.958740234375),
    to_complex(0.281494140625, - 0.959472656250),
    to_complex(0.278564453125, - 0.960449218750),
    to_complex(0.275634765625, - 0.961181640625),
    to_complex(0.272705078125, - 0.962158203125),
    to_complex(0.269775390625, - 0.962890625000),
    to_complex(0.266601562500, - 0.963867187500),
    to_complex(0.263671875000, - 0.964599609375),
    to_complex(0.260742187500, - 0.965332031250),
    to_complex(0.257812500000, - 0.966308593750),
    to_complex(0.254882812500, - 0.967041015625),
    to_complex(0.251953125000, - 0.967773437500),
    to_complex(0.249023437500, - 0.968505859375),
    to_complex(0.245849609375, - 0.969238281250),
    to_complex(0.242919921875, - 0.969970703125),
    to_complex(0.239990234375, - 0.970703125000),
    to_complex(0.237060546875, - 0.971435546875),
    to_complex(0.234130859375, - 0.972167968750),
    to_complex(0.230957031250, - 0.972900390625),
    to_complex(0.228027343750, - 0.973632812500),
    to_complex(0.225097656250, - 0.974365234375),
    to_complex(0.222167968750, - 0.975097656250),
    to_complex(0.218994140625, - 0.975585937500),
    to_complex(0.216064453125, - 0.976318359375),
    to_complex(0.213134765625, - 0.977050781250),
    to_complex(0.210205078125, - 0.977783203125),
    to_complex(0.207031250000, - 0.978271484375),
    to_complex(0.204101562500, - 0.979003906250),
    to_complex(0.201171875000, - 0.979492187500),
    to_complex(0.197998046875, - 0.980224609375),
    to_complex(0.195068359375, - 0.980712890625),
    to_complex(0.192138671875, - 0.981445312500),
    to_complex(0.188964843750, - 0.981933593750),
    to_complex(0.186035156250, - 0.982421875000),
    to_complex(0.183105468750, - 0.983154296875),
    to_complex(0.179931640625, - 0.983642578125),
    to_complex(0.177001953125, - 0.984130859375),
    to_complex(0.174072265625, - 0.984863281250),
    to_complex(0.170898437500, - 0.985351562500),
    to_complex(0.167968750000, - 0.985839843750),
    to_complex(0.164794921875, - 0.986328125000),
    to_complex(0.161865234375, - 0.986816406250),
    to_complex(0.158935546875, - 0.987304687500),
    to_complex(0.155761718750, - 0.987792968750),
    to_complex(0.152832031250, - 0.988281250000),
    to_complex(0.149658203125, - 0.988769531250),
    to_complex(0.146728515625, - 0.989257812500),
    to_complex(0.143798828125, - 0.989501953125),
    to_complex(0.140625000000, - 0.989990234375),
    to_complex(0.137695312500, - 0.990478515625),
    to_complex(0.134521484375, - 0.990966796875),
    to_complex(0.131591796875, - 0.991210937500),
    to_complex(0.128417968750, - 0.991699218750),
    to_complex(0.125488281250, - 0.992187500000),
    to_complex(0.122314453125, - 0.992431640625),
    to_complex(0.119384765625, - 0.992919921875),
    to_complex(0.116210937500, - 0.993164062500),
    to_complex(0.113281250000, - 0.993652343750),
    to_complex(0.110107421875, - 0.993896484375),
    to_complex(0.107177734375, - 0.994140625000),
    to_complex(0.104003906250, - 0.994628906250),
    to_complex(0.101074218750, - 0.994873046875),
    to_complex(0.097900390625, - 0.995117187500),
    to_complex(0.094970703125, - 0.995361328125),
    to_complex(0.091796875000, - 0.995849609375),
    to_complex(0.088867187500, - 0.996093750000),
    to_complex(0.085693359375, - 0.996337890625),
    to_complex(0.082763671875, - 0.996582031250),
    to_complex(0.079589843750, - 0.996826171875),
    to_complex(0.076660156250, - 0.997070312500),
    to_complex(0.073486328125, - 0.997314453125),
    to_complex(0.070556640625, - 0.997558593750),
    to_complex(0.067382812500, - 0.997802734375),
    to_complex(0.064453125000, - 0.998046875000),
    to_complex(0.061279296875, - 0.998046875000),
    to_complex(0.058349609375, - 0.998291015625),
    to_complex(0.055175781250, - 0.998535156250),
    to_complex(0.052246093750, - 0.998535156250),
    to_complex(0.049072265625, - 0.998779296875),
    to_complex(0.045898437500, - 0.999023437500),
    to_complex(0.042968750000, - 0.999023437500),
    to_complex(0.039794921875, - 0.999267578125),
    to_complex(0.036865234375, - 0.999267578125),
    to_complex(0.033691406250, - 0.999511718750),
    to_complex(0.030761718750, - 0.999511718750),
    to_complex(0.027587890625, - 0.999511718750),
    to_complex(0.024658203125, - 0.999755859375),
    to_complex(0.021484375000, - 0.999755859375),
    to_complex(0.018310546875, - 0.999755859375),
    to_complex(0.015380859375, - 1.000000000000),
    to_complex(0.012207031250, - 1.000000000000),
    to_complex(0.009277343750, - 1.000000000000),
    to_complex(0.006103515625, - 1.000000000000),
    to_complex(0.003173828125, - 1.000000000000),
    to_complex(0.000000000000, - 1.000000000000),
    to_complex(- 0.003173828125, - 1.000000000000),
    to_complex(- 0.006103515625, - 1.000000000000),
    to_complex(- 0.009277343750, - 1.000000000000),
    to_complex(- 0.012207031250, - 1.000000000000),
    to_complex(- 0.015380859375, - 1.000000000000),
    to_complex(- 0.018310546875, - 0.999755859375),
    to_complex(- 0.021484375000, - 0.999755859375),
    to_complex(- 0.024658203125, - 0.999755859375),
    to_complex(- 0.027587890625, - 0.999511718750),
    to_complex(- 0.030761718750, - 0.999511718750),
    to_complex(- 0.033691406250, - 0.999511718750),
    to_complex(- 0.036865234375, - 0.999267578125),
    to_complex(- 0.039794921875, - 0.999267578125),
    to_complex(- 0.042968750000, - 0.999023437500),
    to_complex(- 0.045898437500, - 0.999023437500),
    to_complex(- 0.049072265625, - 0.998779296875),
    to_complex(- 0.052246093750, - 0.998535156250),
    to_complex(- 0.055175781250, - 0.998535156250),
    to_complex(- 0.058349609375, - 0.998291015625),
    to_complex(- 0.061279296875, - 0.998046875000),
    to_complex(- 0.064453125000, - 0.998046875000),
    to_complex(- 0.067382812500, - 0.997802734375),
    to_complex(- 0.070556640625, - 0.997558593750),
    to_complex(- 0.073486328125, - 0.997314453125),
    to_complex(- 0.076660156250, - 0.997070312500),
    to_complex(- 0.079589843750, - 0.996826171875),
    to_complex(- 0.082763671875, - 0.996582031250),
    to_complex(- 0.085693359375, - 0.996337890625),
    to_complex(- 0.088867187500, - 0.996093750000),
    to_complex(- 0.091796875000, - 0.995849609375),
    to_complex(- 0.094970703125, - 0.995361328125),
    to_complex(- 0.097900390625, - 0.995117187500),
    to_complex(- 0.101074218750, - 0.994873046875),
    to_complex(- 0.104003906250, - 0.994628906250),
    to_complex(- 0.107177734375, - 0.994140625000),
    to_complex(- 0.110107421875, - 0.993896484375),
    to_complex(- 0.113281250000, - 0.993652343750),
    to_complex(- 0.116210937500, - 0.993164062500),
    to_complex(- 0.119384765625, - 0.992919921875),
    to_complex(- 0.122314453125, - 0.992431640625),
    to_complex(- 0.125488281250, - 0.992187500000),
    to_complex(- 0.128417968750, - 0.991699218750),
    to_complex(- 0.131591796875, - 0.991210937500),
    to_complex(- 0.134521484375, - 0.990966796875),
    to_complex(- 0.137695312500, - 0.990478515625),
    to_complex(- 0.140625000000, - 0.989990234375),
    to_complex(- 0.143798828125, - 0.989501953125),
    to_complex(- 0.146728515625, - 0.989257812500),
    to_complex(- 0.149658203125, - 0.988769531250),
    to_complex(- 0.152832031250, - 0.988281250000),
    to_complex(- 0.155761718750, - 0.987792968750),
    to_complex(- 0.158935546875, - 0.987304687500),
    to_complex(- 0.161865234375, - 0.986816406250),
    to_complex(- 0.164794921875, - 0.986328125000),
    to_complex(- 0.167968750000, - 0.985839843750),
    to_complex(- 0.170898437500, - 0.985351562500),
    to_complex(- 0.174072265625, - 0.984863281250),
    to_complex(- 0.177001953125, - 0.984130859375),
    to_complex(- 0.179931640625, - 0.983642578125),
    to_complex(- 0.183105468750, - 0.983154296875),
    to_complex(- 0.186035156250, - 0.982421875000),
    to_complex(- 0.188964843750, - 0.981933593750),
    to_complex(- 0.192138671875, - 0.981445312500),
    to_complex(- 0.195068359375, - 0.980712890625),
    to_complex(- 0.197998046875, - 0.980224609375),
    to_complex(- 0.201171875000, - 0.979492187500),
    to_complex(- 0.204101562500, - 0.979003906250),
    to_complex(- 0.207031250000, - 0.978271484375),
    to_complex(- 0.210205078125, - 0.977783203125),
    to_complex(- 0.213134765625, - 0.977050781250),
    to_complex(- 0.216064453125, - 0.976318359375),
    to_complex(- 0.218994140625, - 0.975585937500),
    to_complex(- 0.222167968750, - 0.975097656250),
    to_complex(- 0.225097656250, - 0.974365234375),
    to_complex(- 0.228027343750, - 0.973632812500),
    to_complex(- 0.230957031250, - 0.972900390625),
    to_complex(- 0.234130859375, - 0.972167968750),
    to_complex(- 0.237060546875, - 0.971435546875),
    to_complex(- 0.239990234375, - 0.970703125000),
    to_complex(- 0.242919921875, - 0.969970703125),
    to_complex(- 0.245849609375, - 0.969238281250),
    to_complex(- 0.249023437500, - 0.968505859375),
    to_complex(- 0.251953125000, - 0.967773437500),
    to_complex(- 0.254882812500, - 0.967041015625),
    to_complex(- 0.257812500000, - 0.966308593750),
    to_complex(- 0.260742187500, - 0.965332031250),
    to_complex(- 0.263671875000, - 0.964599609375),
    to_complex(- 0.266601562500, - 0.963867187500),
    to_complex(- 0.269775390625, - 0.962890625000),
    to_complex(- 0.272705078125, - 0.962158203125),
    to_complex(- 0.275634765625, - 0.961181640625),
    to_complex(- 0.278564453125, - 0.960449218750),
    to_complex(- 0.281494140625, - 0.959472656250),
    to_complex(- 0.284423828125, - 0.958740234375),
    to_complex(- 0.287353515625, - 0.957763671875),
    to_complex(- 0.290283203125, - 0.957031250000),
    to_complex(- 0.293212890625, - 0.956054687500),
    to_complex(- 0.296142578125, - 0.955078125000),
    to_complex(- 0.299072265625, - 0.954345703125),
    to_complex(- 0.302001953125, - 0.953369140625),
    to_complex(- 0.304931640625, - 0.952392578125),
    to_complex(- 0.307861328125, - 0.951416015625),
    to_complex(- 0.310791015625, - 0.950439453125),
    to_complex(- 0.313720703125, - 0.949462890625),
    to_complex(- 0.316650390625, - 0.948486328125),
    to_complex(- 0.319580078125, - 0.947509765625),
    to_complex(- 0.322509765625, - 0.946533203125),
    to_complex(- 0.325195312500, - 0.945556640625),
    to_complex(- 0.328125000000, - 0.944580078125),
    to_complex(- 0.331054687500, - 0.943603515625),
    to_complex(- 0.333984375000, - 0.942626953125),
    to_complex(- 0.336914062500, - 0.941650390625),
    to_complex(- 0.339843750000, - 0.940429687500),
    to_complex(- 0.342773437500, - 0.939453125000),
    to_complex(- 0.345458984375, - 0.938476562500),
    to_complex(- 0.348388671875, - 0.937255859375),
    to_complex(- 0.351318359375, - 0.936279296875),
    to_complex(- 0.354248046875, - 0.935302734375),
    to_complex(- 0.356933593750, - 0.934082031250),
    to_complex(- 0.359863281250, - 0.933105468750),
    to_complex(- 0.362792968750, - 0.931884765625),
    to_complex(- 0.365722656250, - 0.930664062500),
    to_complex(- 0.368408203125, - 0.929687500000),
    to_complex(- 0.371337890625, - 0.928466796875),
    to_complex(- 0.374267578125, - 0.927246093750),
    to_complex(- 0.376953125000, - 0.926269531250),
    to_complex(- 0.379882812500, - 0.925048828125),
    to_complex(- 0.382568359375, - 0.923828125000),
    to_complex(- 0.385498046875, - 0.922607421875),
    to_complex(- 0.388427734375, - 0.921630859375),
    to_complex(- 0.391113281250, - 0.920410156250),
    to_complex(- 0.394042968750, - 0.919189453125),
    to_complex(- 0.396728515625, - 0.917968750000),
    to_complex(- 0.399658203125, - 0.916748046875),
    to_complex(- 0.402343750000, - 0.915527343750),
    to_complex(- 0.405273437500, - 0.914306640625),
    to_complex(- 0.407958984375, - 0.912841796875),
    to_complex(- 0.410888671875, - 0.911621093750),
    to_complex(- 0.413574218750, - 0.910400390625),
    to_complex(- 0.416503906250, - 0.909179687500),
    to_complex(- 0.419189453125, - 0.907958984375),
    to_complex(- 0.422119140625, - 0.906494140625),
    to_complex(- 0.424804687500, - 0.905273437500),
    to_complex(- 0.427490234375, - 0.904052734375),
    to_complex(- 0.430419921875, - 0.902587890625),
    to_complex(- 0.433105468750, - 0.901367187500),
    to_complex(- 0.435791015625, - 0.899902343750),
    to_complex(- 0.438720703125, - 0.898681640625),
    to_complex(- 0.441406250000, - 0.897216796875),
    to_complex(- 0.444091796875, - 0.895996093750),
    to_complex(- 0.446777343750, - 0.894531250000),
    to_complex(- 0.449707031250, - 0.893310546875),
    to_complex(- 0.452392578125, - 0.891845703125),
    to_complex(- 0.455078125000, - 0.890380859375),
    to_complex(- 0.457763671875, - 0.889160156250),
    to_complex(- 0.460449218750, - 0.887695312500),
    to_complex(- 0.463378906250, - 0.886230468750),
    to_complex(- 0.466064453125, - 0.884765625000),
    to_complex(- 0.468750000000, - 0.883300781250),
    to_complex(- 0.471435546875, - 0.881835937500),
    to_complex(- 0.474121093750, - 0.880371093750),
    to_complex(- 0.476806640625, - 0.878906250000),
    to_complex(- 0.479492187500, - 0.877441406250),
    to_complex(- 0.482177734375, - 0.875976562500),
    to_complex(- 0.484863281250, - 0.874511718750),
    to_complex(- 0.487548828125, - 0.873046875000),
    to_complex(- 0.490234375000, - 0.871582031250),
    to_complex(- 0.492919921875, - 0.870117187500),
    to_complex(- 0.495605468750, - 0.868652343750),
    to_complex(- 0.498291015625, - 0.866943359375),
    to_complex(- 0.500976562500, - 0.865478515625),
    to_complex(- 0.503417968750, - 0.864013671875),
    to_complex(- 0.506103515625, - 0.862304687500),
    to_complex(- 0.508789062500, - 0.860839843750),
    to_complex(- 0.511474609375, - 0.859375000000),
    to_complex(- 0.514160156250, - 0.857666015625),
    to_complex(- 0.516845703125, - 0.856201171875),
    to_complex(- 0.519287109375, - 0.854492187500),
    to_complex(- 0.521972656250, - 0.853027343750),
    to_complex(- 0.524658203125, - 0.851318359375),
    to_complex(- 0.527099609375, - 0.849853515625),
    to_complex(- 0.529785156250, - 0.848144531250),
    to_complex(- 0.532470703125, - 0.846435546875),
    to_complex(- 0.534912109375, - 0.844970703125),
    to_complex(- 0.537597656250, - 0.843261718750),
    to_complex(- 0.540283203125, - 0.841552734375),
    to_complex(- 0.542724609375, - 0.839843750000),
    to_complex(- 0.545410156250, - 0.838134765625),
    to_complex(- 0.547851562500, - 0.836425781250),
    to_complex(- 0.550537109375, - 0.834960937500),
    to_complex(- 0.552978515625, - 0.833251953125),
    to_complex(- 0.555664062500, - 0.831542968750),
    to_complex(- 0.558105468750, - 0.829833984375),
    to_complex(- 0.560546875000, - 0.828125000000),
    to_complex(- 0.563232421875, - 0.826416015625),
    to_complex(- 0.565673828125, - 0.824707031250),
    to_complex(- 0.568359375000, - 0.822753906250),
    to_complex(- 0.570800781250, - 0.821044921875),
    to_complex(- 0.573242187500, - 0.819335937500),
    to_complex(- 0.575927734375, - 0.817626953125),
    to_complex(- 0.578369140625, - 0.815917968750),
    to_complex(- 0.580810546875, - 0.813964843750),
    to_complex(- 0.583251953125, - 0.812255859375),
    to_complex(- 0.585693359375, - 0.810546875000),
    to_complex(- 0.588378906250, - 0.808593750000),
    to_complex(- 0.590820312500, - 0.806884765625),
    to_complex(- 0.593261718750, - 0.804931640625),
    to_complex(- 0.595703125000, - 0.803222656250),
    to_complex(- 0.598144531250, - 0.801269531250),
    to_complex(- 0.600585937500, - 0.799560546875),
    to_complex(- 0.603027343750, - 0.797607421875),
    to_complex(- 0.605468750000, - 0.795898437500),
    to_complex(- 0.607910156250, - 0.793945312500),
    to_complex(- 0.610351562500, - 0.791992187500),
    to_complex(- 0.612792968750, - 0.790283203125),
    to_complex(- 0.615234375000, - 0.788330078125),
    to_complex(- 0.617675781250, - 0.786376953125),
    to_complex(- 0.620117187500, - 0.784667968750),
    to_complex(- 0.622558593750, - 0.782714843750),
    to_complex(- 0.624755859375, - 0.780761718750),
    to_complex(- 0.627197265625, - 0.778808593750),
    to_complex(- 0.629638671875, - 0.776855468750),
    to_complex(- 0.632080078125, - 0.774902343750),
    to_complex(- 0.634277343750, - 0.772949218750),
    to_complex(- 0.636718750000, - 0.770996093750),
    to_complex(- 0.639160156250, - 0.769042968750),
    to_complex(- 0.641601562500, - 0.767089843750),
    to_complex(- 0.643798828125, - 0.765136718750),
    to_complex(- 0.646240234375, - 0.763183593750),
    to_complex(- 0.648437500000, - 0.761230468750),
    to_complex(- 0.650878906250, - 0.759277343750),
    to_complex(- 0.653076171875, - 0.757324218750),
    to_complex(- 0.655517578125, - 0.755126953125),
    to_complex(- 0.657714843750, - 0.753173828125),
    to_complex(- 0.660156250000, - 0.751220703125),
    to_complex(- 0.662353515625, - 0.749023437500),
    to_complex(- 0.664794921875, - 0.747070312500),
    to_complex(- 0.666992187500, - 0.745117187500),
    to_complex(- 0.669189453125, - 0.742919921875),
    to_complex(- 0.671630859375, - 0.740966796875),
    to_complex(- 0.673828125000, - 0.738769531250),
    to_complex(- 0.676025390625, - 0.736816406250),
    to_complex(- 0.678466796875, - 0.734619140625),
    to_complex(- 0.680664062500, - 0.732666015625),
    to_complex(- 0.682861328125, - 0.730468750000),
    to_complex(- 0.685058593750, - 0.728515625000),
    to_complex(- 0.687255859375, - 0.726318359375),
    to_complex(- 0.689453125000, - 0.724365234375),
    to_complex(- 0.691650390625, - 0.722167968750),
    to_complex(- 0.694091796875, - 0.719970703125),
    to_complex(- 0.696289062500, - 0.717773437500),
    to_complex(- 0.698486328125, - 0.715820312500),
    to_complex(- 0.700683593750, - 0.713623046875),
    to_complex(- 0.702636718750, - 0.711425781250),
    to_complex(- 0.704833984375, - 0.709228515625),
    to_complex(- 0.707031250000, - 0.707031250000),
    to_complex(- 0.709228515625, - 0.704833984375),
    to_complex(- 0.711425781250, - 0.702636718750),
    to_complex(- 0.713623046875, - 0.700683593750),
    to_complex(- 0.715820312500, - 0.698486328125),
    to_complex(- 0.717773437500, - 0.696289062500),
    to_complex(- 0.719970703125, - 0.694091796875),
    to_complex(- 0.722167968750, - 0.691650390625),
    to_complex(- 0.724365234375, - 0.689453125000),
    to_complex(- 0.726318359375, - 0.687255859375),
    to_complex(- 0.728515625000, - 0.685058593750),
    to_complex(- 0.730468750000, - 0.682861328125),
    to_complex(- 0.732666015625, - 0.680664062500),
    to_complex(- 0.734619140625, - 0.678466796875),
    to_complex(- 0.736816406250, - 0.676025390625),
    to_complex(- 0.738769531250, - 0.673828125000),
    to_complex(- 0.740966796875, - 0.671630859375),
    to_complex(- 0.742919921875, - 0.669189453125),
    to_complex(- 0.745117187500, - 0.666992187500),
    to_complex(- 0.747070312500, - 0.664794921875),
    to_complex(- 0.749023437500, - 0.662353515625),
    to_complex(- 0.751220703125, - 0.660156250000),
    to_complex(- 0.753173828125, - 0.657714843750),
    to_complex(- 0.755126953125, - 0.655517578125),
    to_complex(- 0.757324218750, - 0.653076171875),
    to_complex(- 0.759277343750, - 0.650878906250),
    to_complex(- 0.761230468750, - 0.648437500000),
    to_complex(- 0.763183593750, - 0.646240234375),
    to_complex(- 0.765136718750, - 0.643798828125),
    to_complex(- 0.767089843750, - 0.641601562500),
    to_complex(- 0.769042968750, - 0.639160156250),
    to_complex(- 0.770996093750, - 0.636718750000),
    to_complex(- 0.772949218750, - 0.634277343750),
    to_complex(- 0.774902343750, - 0.632080078125),
    to_complex(- 0.776855468750, - 0.629638671875),
    to_complex(- 0.778808593750, - 0.627197265625),
    to_complex(- 0.780761718750, - 0.624755859375),
    to_complex(- 0.782714843750, - 0.622558593750),
    to_complex(- 0.784667968750, - 0.620117187500),
    to_complex(- 0.786376953125, - 0.617675781250),
    to_complex(- 0.788330078125, - 0.615234375000),
    to_complex(- 0.790283203125, - 0.612792968750),
    to_complex(- 0.791992187500, - 0.610351562500),
    to_complex(- 0.793945312500, - 0.607910156250),
    to_complex(- 0.795898437500, - 0.605468750000),
    to_complex(- 0.797607421875, - 0.603027343750),
    to_complex(- 0.799560546875, - 0.600585937500),
    to_complex(- 0.801269531250, - 0.598144531250),
    to_complex(- 0.803222656250, - 0.595703125000),
    to_complex(- 0.804931640625, - 0.593261718750),
    to_complex(- 0.806884765625, - 0.590820312500),
    to_complex(- 0.808593750000, - 0.588378906250),
    to_complex(- 0.810546875000, - 0.585693359375),
    to_complex(- 0.812255859375, - 0.583251953125),
    to_complex(- 0.813964843750, - 0.580810546875),
    to_complex(- 0.815917968750, - 0.578369140625),
    to_complex(- 0.817626953125, - 0.575927734375),
    to_complex(- 0.819335937500, - 0.573242187500),
    to_complex(- 0.821044921875, - 0.570800781250),
    to_complex(- 0.822753906250, - 0.568359375000),
    to_complex(- 0.824707031250, - 0.565673828125),
    to_complex(- 0.826416015625, - 0.563232421875),
    to_complex(- 0.828125000000, - 0.560546875000),
    to_complex(- 0.829833984375, - 0.558105468750),
    to_complex(- 0.831542968750, - 0.555664062500),
    to_complex(- 0.833251953125, - 0.552978515625),
    to_complex(- 0.834960937500, - 0.550537109375),
    to_complex(- 0.836425781250, - 0.547851562500),
    to_complex(- 0.838134765625, - 0.545410156250),
    to_complex(- 0.839843750000, - 0.542724609375),
    to_complex(- 0.841552734375, - 0.540283203125),
    to_complex(- 0.843261718750, - 0.537597656250),
    to_complex(- 0.844970703125, - 0.534912109375),
    to_complex(- 0.846435546875, - 0.532470703125),
    to_complex(- 0.848144531250, - 0.529785156250),
    to_complex(- 0.849853515625, - 0.527099609375),
    to_complex(- 0.851318359375, - 0.524658203125),
    to_complex(- 0.853027343750, - 0.521972656250),
    to_complex(- 0.854492187500, - 0.519287109375),
    to_complex(- 0.856201171875, - 0.516845703125),
    to_complex(- 0.857666015625, - 0.514160156250),
    to_complex(- 0.859375000000, - 0.511474609375),
    to_complex(- 0.860839843750, - 0.508789062500),
    to_complex(- 0.862304687500, - 0.506103515625),
    to_complex(- 0.864013671875, - 0.503417968750),
    to_complex(- 0.865478515625, - 0.500976562500),
    to_complex(- 0.866943359375, - 0.498291015625),
    to_complex(- 0.868652343750, - 0.495605468750),
    to_complex(- 0.870117187500, - 0.492919921875),
    to_complex(- 0.871582031250, - 0.490234375000),
    to_complex(- 0.873046875000, - 0.487548828125),
    to_complex(- 0.874511718750, - 0.484863281250),
    to_complex(- 0.875976562500, - 0.482177734375),
    to_complex(- 0.877441406250, - 0.479492187500),
    to_complex(- 0.878906250000, - 0.476806640625),
    to_complex(- 0.880371093750, - 0.474121093750),
    to_complex(- 0.881835937500, - 0.471435546875),
    to_complex(- 0.883300781250, - 0.468750000000),
    to_complex(- 0.884765625000, - 0.466064453125),
    to_complex(- 0.886230468750, - 0.463378906250),
    to_complex(- 0.887695312500, - 0.460449218750),
    to_complex(- 0.889160156250, - 0.457763671875),
    to_complex(- 0.890380859375, - 0.455078125000),
    to_complex(- 0.891845703125, - 0.452392578125),
    to_complex(- 0.893310546875, - 0.449707031250),
    to_complex(- 0.894531250000, - 0.446777343750),
    to_complex(- 0.895996093750, - 0.444091796875),
    to_complex(- 0.897216796875, - 0.441406250000),
    to_complex(- 0.898681640625, - 0.438720703125),
    to_complex(- 0.899902343750, - 0.435791015625),
    to_complex(- 0.901367187500, - 0.433105468750),
    to_complex(- 0.902587890625, - 0.430419921875),
    to_complex(- 0.904052734375, - 0.427490234375),
    to_complex(- 0.905273437500, - 0.424804687500),
    to_complex(- 0.906494140625, - 0.422119140625),
    to_complex(- 0.907958984375, - 0.419189453125),
    to_complex(- 0.909179687500, - 0.416503906250),
    to_complex(- 0.910400390625, - 0.413574218750),
    to_complex(- 0.911621093750, - 0.410888671875),
    to_complex(- 0.912841796875, - 0.407958984375),
    to_complex(- 0.914306640625, - 0.405273437500),
    to_complex(- 0.915527343750, - 0.402343750000),
    to_complex(- 0.916748046875, - 0.399658203125),
    to_complex(- 0.917968750000, - 0.396728515625),
    to_complex(- 0.919189453125, - 0.394042968750),
    to_complex(- 0.920410156250, - 0.391113281250),
    to_complex(- 0.921630859375, - 0.388427734375),
    to_complex(- 0.922607421875, - 0.385498046875),
    to_complex(- 0.923828125000, - 0.382568359375),
    to_complex(- 0.925048828125, - 0.379882812500),
    to_complex(- 0.926269531250, - 0.376953125000),
    to_complex(- 0.927246093750, - 0.374267578125),
    to_complex(- 0.928466796875, - 0.371337890625),
    to_complex(- 0.929687500000, - 0.368408203125),
    to_complex(- 0.930664062500, - 0.365722656250),
    to_complex(- 0.931884765625, - 0.362792968750),
    to_complex(- 0.933105468750, - 0.359863281250),
    to_complex(- 0.934082031250, - 0.356933593750),
    to_complex(- 0.935302734375, - 0.354248046875),
    to_complex(- 0.936279296875, - 0.351318359375),
    to_complex(- 0.937255859375, - 0.348388671875),
    to_complex(- 0.938476562500, - 0.345458984375),
    to_complex(- 0.939453125000, - 0.342773437500),
    to_complex(- 0.940429687500, - 0.339843750000),
    to_complex(- 0.941650390625, - 0.336914062500),
    to_complex(- 0.942626953125, - 0.333984375000),
    to_complex(- 0.943603515625, - 0.331054687500),
    to_complex(- 0.944580078125, - 0.328125000000),
    to_complex(- 0.945556640625, - 0.325195312500),
    to_complex(- 0.946533203125, - 0.322509765625),
    to_complex(- 0.947509765625, - 0.319580078125),
    to_complex(- 0.948486328125, - 0.316650390625),
    to_complex(- 0.949462890625, - 0.313720703125),
    to_complex(- 0.950439453125, - 0.310791015625),
    to_complex(- 0.951416015625, - 0.307861328125),
    to_complex(- 0.952392578125, - 0.304931640625),
    to_complex(- 0.953369140625, - 0.302001953125),
    to_complex(- 0.954345703125, - 0.299072265625),
    to_complex(- 0.955078125000, - 0.296142578125),
    to_complex(- 0.956054687500, - 0.293212890625),
    to_complex(- 0.957031250000, - 0.290283203125),
    to_complex(- 0.957763671875, - 0.287353515625),
    to_complex(- 0.958740234375, - 0.284423828125),
    to_complex(- 0.959472656250, - 0.281494140625),
    to_complex(- 0.960449218750, - 0.278564453125),
    to_complex(- 0.961181640625, - 0.275634765625),
    to_complex(- 0.962158203125, - 0.272705078125),
    to_complex(- 0.962890625000, - 0.269775390625),
    to_complex(- 0.963867187500, - 0.266601562500),
    to_complex(- 0.964599609375, - 0.263671875000),
    to_complex(- 0.965332031250, - 0.260742187500),
    to_complex(- 0.966308593750, - 0.257812500000),
    to_complex(- 0.967041015625, - 0.254882812500),
    to_complex(- 0.967773437500, - 0.251953125000),
    to_complex(- 0.968505859375, - 0.249023437500),
    to_complex(- 0.969238281250, - 0.245849609375),
    to_complex(- 0.969970703125, - 0.242919921875),
    to_complex(- 0.970703125000, - 0.239990234375),
    to_complex(- 0.971435546875, - 0.237060546875),
    to_complex(- 0.972167968750, - 0.234130859375),
    to_complex(- 0.972900390625, - 0.230957031250),
    to_complex(- 0.973632812500, - 0.228027343750),
    to_complex(- 0.974365234375, - 0.225097656250),
    to_complex(- 0.975097656250, - 0.222167968750),
    to_complex(- 0.975585937500, - 0.218994140625),
    to_complex(- 0.976318359375, - 0.216064453125),
    to_complex(- 0.977050781250, - 0.213134765625),
    to_complex(- 0.977783203125, - 0.210205078125),
    to_complex(- 0.978271484375, - 0.207031250000),
    to_complex(- 0.979003906250, - 0.204101562500),
    to_complex(- 0.979492187500, - 0.201171875000),
    to_complex(- 0.980224609375, - 0.197998046875),
    to_complex(- 0.980712890625, - 0.195068359375),
    to_complex(- 0.981445312500, - 0.192138671875),
    to_complex(- 0.981933593750, - 0.188964843750),
    to_complex(- 0.982421875000, - 0.186035156250),
    to_complex(- 0.983154296875, - 0.183105468750),
    to_complex(- 0.983642578125, - 0.179931640625),
    to_complex(- 0.984130859375, - 0.177001953125),
    to_complex(- 0.984863281250, - 0.174072265625),
    to_complex(- 0.985351562500, - 0.170898437500),
    to_complex(- 0.985839843750, - 0.167968750000),
    to_complex(- 0.986328125000, - 0.164794921875),
    to_complex(- 0.986816406250, - 0.161865234375),
    to_complex(- 0.987304687500, - 0.158935546875),
    to_complex(- 0.987792968750, - 0.155761718750),
    to_complex(- 0.988281250000, - 0.152832031250),
    to_complex(- 0.988769531250, - 0.149658203125),
    to_complex(- 0.989257812500, - 0.146728515625),
    to_complex(- 0.989501953125, - 0.143798828125),
    to_complex(- 0.989990234375, - 0.140625000000),
    to_complex(- 0.990478515625, - 0.137695312500),
    to_complex(- 0.990966796875, - 0.134521484375),
    to_complex(- 0.991210937500, - 0.131591796875),
    to_complex(- 0.991699218750, - 0.128417968750),
    to_complex(- 0.992187500000, - 0.125488281250),
    to_complex(- 0.992431640625, - 0.122314453125),
    to_complex(- 0.992919921875, - 0.119384765625),
    to_complex(- 0.993164062500, - 0.116210937500),
    to_complex(- 0.993652343750, - 0.113281250000),
    to_complex(- 0.993896484375, - 0.110107421875),
    to_complex(- 0.994140625000, - 0.107177734375),
    to_complex(- 0.994628906250, - 0.104003906250),
    to_complex(- 0.994873046875, - 0.101074218750),
    to_complex(- 0.995117187500, - 0.097900390625),
    to_complex(- 0.995361328125, - 0.094970703125),
    to_complex(- 0.995849609375, - 0.091796875000),
    to_complex(- 0.996093750000, - 0.088867187500),
    to_complex(- 0.996337890625, - 0.085693359375),
    to_complex(- 0.996582031250, - 0.082763671875),
    to_complex(- 0.996826171875, - 0.079589843750),
    to_complex(- 0.997070312500, - 0.076660156250),
    to_complex(- 0.997314453125, - 0.073486328125),
    to_complex(- 0.997558593750, - 0.070556640625),
    to_complex(- 0.997802734375, - 0.067382812500),
    to_complex(- 0.998046875000, - 0.064453125000),
    to_complex(- 0.998046875000, - 0.061279296875),
    to_complex(- 0.998291015625, - 0.058349609375),
    to_complex(- 0.998535156250, - 0.055175781250),
    to_complex(- 0.998535156250, - 0.052246093750),
    to_complex(- 0.998779296875, - 0.049072265625),
    to_complex(- 0.999023437500, - 0.045898437500),
    to_complex(- 0.999023437500, - 0.042968750000),
    to_complex(- 0.999267578125, - 0.039794921875),
    to_complex(- 0.999267578125, - 0.036865234375),
    to_complex(- 0.999511718750, - 0.033691406250),
    to_complex(- 0.999511718750, - 0.030761718750),
    to_complex(- 0.999511718750, - 0.027587890625),
    to_complex(- 0.999755859375, - 0.024658203125),
    to_complex(- 0.999755859375, - 0.021484375000),
    to_complex(- 0.999755859375, - 0.018310546875),
    to_complex(- 1.000000000000, - 0.015380859375),
    to_complex(- 1.000000000000, - 0.012207031250),
    to_complex(- 1.000000000000, - 0.009277343750),
    to_complex(- 1.000000000000, - 0.006103515625),
    to_complex(- 1.000000000000, - 0.003173828125));

end package;