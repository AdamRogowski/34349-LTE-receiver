library IEEE;
  use work.complex_pkg.all;

package test_constants is

  constant TWIDDLE_VALUES_4 : complex_array(0 to 1) := (
to_complex(1.000000000000, 0.000000000000) ,
 to_complex(0.000000000000, -1.000000000000));

  constant INPUT_4_16qam_clear : complex_array(0 to 3) := (
to_complex(0.000000000000, 0.000000000000) ,
 to_complex(1.000000000000, 0.000000000000) ,
 to_complex(2.000000000000, 2.000000000000) ,
 to_complex(0.000000000000, 1.000000000000));

  constant TWIDDLE_VALUES_64 : complex_array(0 to 63) := (
    to_complex(1.000000000000, 0.000000000000),
    to_complex(0.995117187500, - 0.097900390625),
    to_complex(0.980712890625, - 0.195068359375),
    to_complex(0.957031250000, - 0.290283203125),
    to_complex(0.923828125000, - 0.382568359375),
    to_complex(0.881835937500, - 0.471435546875),
    to_complex(0.831542968750, - 0.555664062500),
    to_complex(0.772949218750, - 0.634277343750),
    to_complex(0.707031250000, - 0.707031250000),
    to_complex(0.634277343750, - 0.772949218750),
    to_complex(0.555664062500, - 0.831542968750),
    to_complex(0.471435546875, - 0.881835937500),
    to_complex(0.382568359375, - 0.923828125000),
    to_complex(0.290283203125, - 0.957031250000),
    to_complex(0.195068359375, - 0.980712890625),
    to_complex(0.097900390625, - 0.995117187500),
    to_complex(0.000000000000, - 1.000000000000),
    to_complex(- 0.097900390625, - 0.995117187500),
    to_complex(- 0.195068359375, - 0.980712890625),
    to_complex(- 0.290283203125, - 0.957031250000),
    to_complex(- 0.382568359375, - 0.923828125000),
    to_complex(- 0.471435546875, - 0.881835937500),
    to_complex(- 0.555664062500, - 0.831542968750),
    to_complex(- 0.634277343750, - 0.772949218750),
    to_complex(- 0.707031250000, - 0.707031250000),
    to_complex(- 0.772949218750, - 0.634277343750),
    to_complex(- 0.831542968750, - 0.555664062500),
    to_complex(- 0.881835937500, - 0.471435546875),
    to_complex(- 0.923828125000, - 0.382568359375),
    to_complex(- 0.957031250000, - 0.290283203125),
    to_complex(- 0.980712890625, - 0.195068359375),
    to_complex(- 0.995117187500, - 0.097900390625),
    to_complex(- 1.000000000000, 0.000000000000),
    to_complex(- 0.995117187500, 0.097900390625),
    to_complex(- 0.980712890625, 0.195068359375),
    to_complex(- 0.957031250000, 0.290283203125),
    to_complex(- 0.923828125000, 0.382568359375),
    to_complex(- 0.881835937500, 0.471435546875),
    to_complex(- 0.831542968750, 0.555664062500),
    to_complex(- 0.772949218750, 0.634277343750),
    to_complex(- 0.707031250000, 0.707031250000),
    to_complex(- 0.634277343750, 0.772949218750),
    to_complex(- 0.555664062500, 0.831542968750),
    to_complex(- 0.471435546875, 0.881835937500),
    to_complex(- 0.382568359375, 0.923828125000),
    to_complex(- 0.290283203125, 0.957031250000),
    to_complex(- 0.195068359375, 0.980712890625),
    to_complex(- 0.097900390625, 0.995117187500),
    to_complex(0.000000000000, 1.000000000000),
    to_complex(0.097900390625, 0.995117187500),
    to_complex(0.195068359375, 0.980712890625),
    to_complex(0.290283203125, 0.957031250000),
    to_complex(0.382568359375, 0.923828125000),
    to_complex(0.471435546875, 0.881835937500),
    to_complex(0.555664062500, 0.831542968750),
    to_complex(0.634277343750, 0.772949218750),
    to_complex(0.707031250000, 0.707031250000),
    to_complex(0.772949218750, 0.634277343750),
    to_complex(0.831542968750, 0.555664062500),
    to_complex(0.881835937500, 0.471435546875),
    to_complex(0.923828125000, 0.382568359375),
    to_complex(0.957031250000, 0.290283203125),
    to_complex(0.980712890625, 0.195068359375),
    to_complex(0.995117187500, 0.097900390625));

  -- input_bits = [0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 0 1 0 1 0 1 0 1 0 1 0 1 0 1 0 1 0 1 0 1 0 1 0 1 0 1 0 1 0 1 0 1 1 0 1 0 1 0 1 0 1 0 1 0 1 0 1 0 1 0 1 0 1 0 1 0 1 0 1 0 1 0 1 0];
  constant INPUT_64_qpsk : complex_array(0 to 63) := (
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.449707031250, - 0.022216796875),
    to_complex(- 0.448730468750, 0.044189453125),
    to_complex(- 0.148925781250, 0.022216796875),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.088134765625, - 0.022216796875),
    to_complex(- 0.145751953125, 0.044189453125),
    to_complex(- 0.061767578125, 0.022216796875),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.046630859375, - 0.022216796875),
    to_complex(- 0.082763671875, 0.044189453125),
    to_complex(- 0.036865234375, 0.022216796875),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.029785156250, - 0.022216796875),
    to_complex(- 0.053955078125, 0.044189453125),
    to_complex(- 0.024414062500, 0.022216796875),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.020019531250, - 0.022216796875),
    to_complex(- 0.036376953125, 0.044189453125),
    to_complex(- 0.016357421875, 0.022216796875),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.013183593750, - 0.022216796875),
    to_complex(- 0.023681640625, 0.044189453125),
    to_complex(- 0.010498046875, 0.022216796875),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.007812500000, - 0.022216796875),
    to_complex(- 0.013427734375, 0.044189453125),
    to_complex(- 0.005615234375, 0.022216796875),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.003173828125, - 0.022216796875),
    to_complex(- 0.004394531250, 0.044189453125),
    to_complex(- 0.000976562500, 0.022216796875),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.000976562500, - 0.022216796875),
    to_complex(0.004394531250, 0.044189453125),
    to_complex(0.003173828125, 0.022216796875),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.005615234375, - 0.022216796875),
    to_complex(0.013427734375, 0.044189453125),
    to_complex(0.007812500000, 0.022216796875),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.010498046875, - 0.022216796875),
    to_complex(0.023681640625, 0.044189453125),
    to_complex(0.013183593750, 0.022216796875),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.016357421875, - 0.022216796875),
    to_complex(0.036376953125, 0.044189453125),
    to_complex(0.020019531250, 0.022216796875),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.024414062500, - 0.022216796875),
    to_complex(0.053955078125, 0.044189453125),
    to_complex(0.029785156250, 0.022216796875),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.036865234375, - 0.022216796875),
    to_complex(0.082763671875, 0.044189453125),
    to_complex(0.046630859375, 0.022216796875),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.061767578125, - 0.022216796875),
    to_complex(0.145751953125, 0.044189453125),
    to_complex(0.088134765625, 0.022216796875),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.148925781250, - 0.022216796875),
    to_complex(0.448730468750, 0.044189453125),
    to_complex(0.449707031250, 0.022216796875));

  constant INPUT_64_16qam_clear : complex_array(0 to 63) := (--without noise
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.667358363281, 0.604858363281),
    to_complex(- 1.144146298451, 1.394146298451),
    to_complex(- 0.241920387669, - 0.179420387669),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.156006993243, 0.093506993243),
    to_complex(- 0.287069776117, 0.537069776117),
    to_complex(- 0.118587899140, - 0.056087899140),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.097322573673, 0.034822573673),
    to_complex(- 0.108858551474, 0.358858551474),
    to_complex(- 0.083387475174, - 0.020887475174),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.073385747296, 0.010885747296),
    to_complex(- 0.027312940698, 0.277312940698),
    to_complex(- 0.065729061742, - 0.003229061742),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.059573349032, - 0.002926650968),
    to_complex(0.022415151146, 0.227584848854),
    to_complex(- 0.054426579571, 0.008073420429),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.049980529178, - 0.012519470822),
    to_complex(0.058186108006, 0.191813891994),
    to_complex(- 0.046030149247, 0.016469850753),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.042431428791, - 0.020068571209),
    to_complex(0.087081664549, 0.162918335451),
    to_complex(- 0.039077717506, 0.023422282494),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.035885499611, - 0.026614500389),
    to_complex(0.112688574580, 0.137311425420),
    to_complex(- 0.032785214055, 0.029714785945),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.029714785945, - 0.032785214055),
    to_complex(0.137311425420, 0.112688574580),
    to_complex(- 0.026614500389, 0.035885499611),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.023422282494, - 0.039077717506),
    to_complex(0.162918335451, 0.087081664549),
    to_complex(- 0.020068571209, 0.042431428791),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.016469850753, - 0.046030149247),
    to_complex(0.191813891994, 0.058186108006),
    to_complex(- 0.012519470822, 0.049980529178),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(0.008073420429, - 0.054426579571),
    to_complex(0.227584848854, 0.022415151146),
    to_complex(- 0.002926650968, 0.059573349032),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.003229061742, - 0.065729061742),
    to_complex(0.277312940698, - 0.027312940698),
    to_complex(0.010885747296, 0.073385747296),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.020887475174, - 0.083387475174),
    to_complex(0.358858551474, - 0.108858551474),
    to_complex(0.034822573673, 0.097322573673),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.056087899140, - 0.118587899140),
    to_complex(0.537069776117, - 0.287069776117),
    to_complex(0.093506993243, 0.156006993243),
    to_complex(0.000000000000, 0.000000000000),
    to_complex(- 0.179420387669, - 0.241920387669),
    to_complex(1.394146298451, - 1.144146298451),
    to_complex(0.604858363281, 0.667358363281));

  constant INPUT_64_16qam_noise : complex_array(0 to 63) := (
to_complex(0.080469106309, -0.040357748519) ,
 to_complex(0.577558222884, 0.586126957643) ,
 to_complex(-1.055495653899, 1.399594892027) ,
 to_complex(-0.228497661160, -0.191025907646) ,
 to_complex(0.039765954840, 0.012001373120) ,
 to_complex(0.089833928502, 0.109409661866) ,
 to_complex(-0.310531637011, 0.500091215782) ,
 to_complex(-0.129644713648, -0.063119295863) ,
 to_complex(0.016808670791, -0.084779621284) ,
 to_complex(0.030909487365, 0.080366205785) ,
 to_complex(-0.090104702750, 0.333843678076) ,
 to_complex(-0.131614568993, -0.068756807482) ,
 to_complex(0.002631950402, -0.010097738673) ,
 to_complex(0.099325724446, -0.045922304363) ,
 to_complex(-0.014307879776, 0.276483568057) ,
 to_complex(-0.022679724947, -0.025523084761) ,
 to_complex(0.040005183856, 0.086596183057) ,
 to_complex(0.033690955530, 0.042342758945) ,
 to_complex(0.032636613029, 0.128299811402) ,
 to_complex(-0.091978380888, 0.025622139960) ,
 to_complex(-0.052558986034, -0.055594906371) ,
 to_complex(0.086754878883, -0.022661366761) ,
 to_complex(0.058188090182, 0.198351179354) ,
 to_complex(-0.048213919509, 0.046202400054) ,
 to_complex(0.036229642228, -0.010857312322) ,
 to_complex(0.066074179309, 0.042610697106) ,
 to_complex(0.101006901687, 0.143794573492) ,
 to_complex(0.010636692768, 0.036445322645) ,
 to_complex(0.036971717015, 0.026432179427) ,
 to_complex(0.045419334619, -0.023227100679) ,
 to_complex(0.085237375701, 0.172341223602) ,
 to_complex(-0.058693291031, 0.042566883329) ,
 to_complex(0.047402186167, -0.031180425347) ,
 to_complex(-0.034377290448, -0.104573243098) ,
 to_complex(0.136338732311, 0.186592803014) ,
 to_complex(-0.104107556121, 0.011847245398) ,
 to_complex(0.040578609983, 0.004109948084) ,
 to_complex(0.057687170084, -0.016684207764) ,
 to_complex(0.162964544000, 0.091598682868) ,
 to_complex(-0.022885309316, 0.006456315062) ,
 to_complex(-0.098863441277, -0.018597985842) ,
 to_complex(0.039579317583, -0.050996215214) ,
 to_complex(0.104634926165, 0.116994727874) ,
 to_complex(-0.104742257806, 0.015751453121) ,
 to_complex(0.003178447002, 0.031201193191) ,
 to_complex(-0.029641537722, -0.042154632100) ,
 to_complex(0.243947171173, 0.013116048840) ,
 to_complex(0.023992380676, 0.017544374734) ,
 to_complex(0.034106479316, -0.011298449203) ,
 to_complex(-0.030711992809, -0.069176173947) ,
 to_complex(0.295181784192, -0.085741285285) ,
 to_complex(0.014887285189, 0.081027592993) ,
 to_complex(0.032847464485, -0.032697288655) ,
 to_complex(0.000432026410, -0.087134814228) ,
 to_complex(0.394561770618, -0.095489520040) ,
 to_complex(0.029576257455, 0.061350329024) ,
 to_complex(-0.005853250465, -0.011462092322) ,
 to_complex(-0.016015264617, -0.104668165925) ,
 to_complex(0.452625724755, -0.360070028026) ,
 to_complex(0.073442853321, 0.197201059020) ,
 to_complex(-0.050523328703, 0.096405149080) ,
 to_complex(-0.194633312412, -0.203771230554) ,
 to_complex(1.419940079924, -1.156702509681) ,
 to_complex(0.637692194868, 0.684401916830));

end package;

